library ieee;
use ieee.std_logic_1164.all;


package mux_pkg is
type array2d is array (natural range <>) of std_logic_vector;
	
end package mux_pkg;

package body mux_pkg is
	
end package body mux_pkg;
