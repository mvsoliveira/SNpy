library ieee;
use ieee.std_logic_1164.all;
use IEEE.math_real.all;

package csn_pkg is

	constant MUON_NUMBER : integer := 352;
	constant IDX_WIDTH   : integer := integer(ceil(log(real(MUON_NUMBER), real(2))));
	constant PT_WIDTH    : integer := 4;
	constant word_w      : integer := PT_WIDTH + IDX_WIDTH;

	type muon_type is record
		idx : std_logic_vector(IDX_WIDTH - 1 downto 0);
		pt  : std_logic_vector(PT_WIDTH - 1 downto 0);
	end record;
	
	type muon_sel_type is record		
		pt  : std_logic_vector(PT_WIDTH - 1 downto 0);
	end record;

	type muon_a is array (natural range <>) of muon_type;
	type muon_sel_a is array (natural range <>) of muon_sel_type;

	type cmp_cfg is record
		a : natural;
		b : natural;
		p : boolean;
	end record;

	-- has to be array of array instead of (x,y) array because of issues with synplify
	type pair_cmp_cfg is array (natural range <>) of cmp_cfg;
	type cfg_net_t is array (natural range <>) of pair_cmp_cfg;
	type stages_a is array(natural range <>) of boolean;

	
	function to_array(data : std_logic_vector; N : integer) return muon_a;    
    function to_sel_array(data : std_logic_vector; N : integer) return muon_sel_a;
    function to_stdv(muon : muon_a; N : integer) return std_logic_vector;
	
	

	--type cfg_net_t is array (natural range <>, natural range <>) of cmp_cfg;
	function get_cfg(I : integer) return cfg_net_t;
	function get_stg(I : integer; D: integer) return stages_a;


	constant empty_cfg : cfg_net_t := (
		((a => 0, b => 1, p => False), (a => 2, b => 3, p => False)),
		((a => 0, b => 2, p => False), (a => 1, b => 3, p => False)),
		((a => 1, b => 2, p => False), (a => 0, b => 3, p => True))
	);

end package csn_pkg;

package body csn_pkg is

	function get_cfg(I : integer) return cfg_net_t is
	begin
		case I is			

			when 64 => return (
                    ((a => 0  , b => 1  , p => False), (a => 2  , b => 3  , p => False), (a => 4  , b => 5  , p => False), (a => 6  , b => 7  , p => False), (a => 8  , b => 9  , p => False), (a => 10 , b => 11 , p => False), (a => 12 , b => 13 , p => False), (a => 14 , b => 15 , p => False), (a => 16 , b => 17 , p => False), (a => 18 , b => 19 , p => False), (a => 20 , b => 21 , p => False), (a => 22 , b => 23 , p => False), (a => 24 , b => 25 , p => False), (a => 26 , b => 27 , p => False), (a => 28 , b => 29 , p => False), (a => 30 , b => 31 , p => False), (a => 32 , b => 33 , p => False), (a => 34 , b => 35 , p => False), (a => 36 , b => 37 , p => False), (a => 38 , b => 39 , p => False), (a => 40 , b => 41 , p => False), (a => 42 , b => 43 , p => False), (a => 44 , b => 45 , p => False), (a => 46 , b => 47 , p => False), (a => 48 , b => 49 , p => False), (a => 50 , b => 51 , p => False), (a => 52 , b => 53 , p => False), (a => 54 , b => 55 , p => False), (a => 56 , b => 57 , p => False), (a => 58 , b => 59 , p => False), (a => 60 , b => 61 , p => False), (a => 62 , b => 63 , p => False)),
                    ((a => 0  , b => 2  , p => False), (a => 4  , b => 6  , p => False), (a => 8  , b => 10 , p => False), (a => 12 , b => 14 , p => False), (a => 16 , b => 18 , p => False), (a => 20 , b => 22 , p => False), (a => 24 , b => 26 , p => False), (a => 28 , b => 30 , p => False), (a => 32 , b => 34 , p => False), (a => 36 , b => 38 , p => False), (a => 40 , b => 42 , p => False), (a => 44 , b => 46 , p => False), (a => 48 , b => 50 , p => False), (a => 52 , b => 54 , p => False), (a => 56 , b => 58 , p => False), (a => 60 , b => 62 , p => False), (a => 1  , b => 3  , p => False), (a => 5  , b => 7  , p => False), (a => 9  , b => 11 , p => False), (a => 13 , b => 15 , p => False), (a => 17 , b => 19 , p => False), (a => 21 , b => 23 , p => False), (a => 25 , b => 27 , p => False), (a => 29 , b => 31 , p => False), (a => 33 , b => 35 , p => False), (a => 37 , b => 39 , p => False), (a => 41 , b => 43 , p => False), (a => 45 , b => 47 , p => False), (a => 49 , b => 51 , p => False), (a => 53 , b => 55 , p => False), (a => 57 , b => 59 , p => False), (a => 61 , b => 63 , p => False)),
                    ((a => 1  , b => 2  , p => False), (a => 5  , b => 6  , p => False), (a => 9  , b => 10 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 21 , b => 22 , p => False), (a => 25 , b => 26 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 37 , b => 38 , p => False), (a => 41 , b => 42 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 53 , b => 54 , p => False), (a => 57 , b => 58 , p => False), (a => 61 , b => 62 , p => False), (a => 0  , b => 4  , p => False), (a => 8  , b => 12 , p => False), (a => 16 , b => 20 , p => False), (a => 24 , b => 28 , p => False), (a => 32 , b => 36 , p => False), (a => 40 , b => 44 , p => False), (a => 48 , b => 52 , p => False), (a => 56 , b => 60 , p => False), (a => 3  , b => 7  , p => False), (a => 11 , b => 15 , p => False), (a => 19 , b => 23 , p => False), (a => 27 , b => 31 , p => False), (a => 35 , b => 39 , p => False), (a => 43 , b => 47 , p => False), (a => 51 , b => 55 , p => False), (a => 59 , b => 63 , p => False)),
                    ((a => 2  , b => 6  , p => False), (a => 10 , b => 14 , p => False), (a => 18 , b => 22 , p => False), (a => 26 , b => 30 , p => False), (a => 34 , b => 38 , p => False), (a => 42 , b => 46 , p => False), (a => 50 , b => 54 , p => False), (a => 58 , b => 62 , p => False), (a => 1  , b => 5  , p => False), (a => 9  , b => 13 , p => False), (a => 17 , b => 21 , p => False), (a => 25 , b => 29 , p => False), (a => 33 , b => 37 , p => False), (a => 41 , b => 45 , p => False), (a => 49 , b => 53 , p => False), (a => 57 , b => 61 , p => False), (a => 0  , b => 8  , p => False), (a => 16 , b => 24 , p => False), (a => 32 , b => 40 , p => False), (a => 48 , b => 56 , p => False), (a => 7  , b => 15 , p => False), (a => 23 , b => 31 , p => False), (a => 39 , b => 47 , p => False), (a => 55 , b => 63 , p => False), (a => 3  , b => 60 , p => True ), (a => 4  , b => 59 , p => True ), (a => 11 , b => 52 , p => True ), (a => 12 , b => 51 , p => True ), (a => 19 , b => 44 , p => True ), (a => 20 , b => 43 , p => True ), (a => 27 , b => 36 , p => True ), (a => 28 , b => 35 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 10 , b => 12 , p => False), (a => 18 , b => 20 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 42 , b => 44 , p => False), (a => 50 , b => 52 , p => False), (a => 58 , b => 60 , p => False), (a => 3  , b => 5  , p => False), (a => 11 , b => 13 , p => False), (a => 19 , b => 21 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 43 , b => 45 , p => False), (a => 51 , b => 53 , p => False), (a => 59 , b => 61 , p => False), (a => 0  , b => 16 , p => False), (a => 32 , b => 48 , p => False), (a => 15 , b => 31 , p => False), (a => 47 , b => 63 , p => False), (a => 1  , b => 62 , p => True ), (a => 6  , b => 57 , p => True ), (a => 7  , b => 56 , p => True ), (a => 8  , b => 55 , p => True ), (a => 9  , b => 54 , p => True ), (a => 14 , b => 49 , p => True ), (a => 17 , b => 46 , p => True ), (a => 22 , b => 41 , p => True ), (a => 23 , b => 40 , p => True ), (a => 24 , b => 39 , p => True ), (a => 25 , b => 38 , p => True ), (a => 30 , b => 33 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 0  , b => 32 , p => False), (a => 7  , b => 63 , p => True ), (a => 8  , b => 56 , p => True ), (a => 15 , b => 55 , p => True ), (a => 16 , b => 48 , p => True ), (a => 23 , b => 47 , p => True ), (a => 24 , b => 40 , p => True ), (a => 31 , b => 39 , p => True )),
                    ((a => 4  , b => 12 , p => False), (a => 20 , b => 28 , p => False), (a => 36 , b => 44 , p => False), (a => 52 , b => 60 , p => False), (a => 2  , b => 10 , p => False), (a => 18 , b => 26 , p => False), (a => 34 , b => 42 , p => False), (a => 50 , b => 58 , p => False), (a => 6  , b => 14 , p => False), (a => 22 , b => 30 , p => False), (a => 38 , b => 46 , p => False), (a => 54 , b => 62 , p => False), (a => 1  , b => 9  , p => False), (a => 17 , b => 25 , p => False), (a => 33 , b => 41 , p => False), (a => 49 , b => 57 , p => False), (a => 5  , b => 13 , p => False), (a => 21 , b => 29 , p => False), (a => 37 , b => 45 , p => False), (a => 53 , b => 61 , p => False), (a => 3  , b => 11 , p => False), (a => 19 , b => 27 , p => False), (a => 35 , b => 43 , p => False), (a => 51 , b => 59 , p => False), (a => 0  , b => 63 , p => True ), (a => 7  , b => 56 , p => True ), (a => 8  , b => 55 , p => True ), (a => 15 , b => 48 , p => True ), (a => 16 , b => 47 , p => True ), (a => 23 , b => 40 , p => True ), (a => 24 , b => 39 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 20 , b => 24 , p => False), (a => 36 , b => 40 , p => False), (a => 52 , b => 56 , p => False), (a => 6  , b => 10 , p => False), (a => 22 , b => 26 , p => False), (a => 38 , b => 42 , p => False), (a => 54 , b => 58 , p => False), (a => 5  , b => 9  , p => False), (a => 21 , b => 25 , p => False), (a => 37 , b => 41 , p => False), (a => 53 , b => 57 , p => False), (a => 7  , b => 11 , p => False), (a => 23 , b => 27 , p => False), (a => 39 , b => 43 , p => False), (a => 55 , b => 59 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 2  , b => 61 , p => True ), (a => 3  , b => 60 , p => True ), (a => 12 , b => 51 , p => True ), (a => 13 , b => 50 , p => True ), (a => 14 , b => 49 , p => True ), (a => 15 , b => 48 , p => True ), (a => 16 , b => 47 , p => True ), (a => 17 , b => 46 , p => True ), (a => 18 , b => 45 , p => True ), (a => 19 , b => 44 , p => True ), (a => 28 , b => 35 , p => True ), (a => 29 , b => 34 , p => True ), (a => 30 , b => 33 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 14 , b => 49 , p => True ), (a => 15 , b => 48 , p => True ), (a => 16 , b => 47 , p => True ), (a => 17 , b => 46 , p => True ), (a => 30 , b => 33 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 0  , b => 63 , p => True ), (a => 15 , b => 48 , p => True ), (a => 16 , b => 47 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 8  , b => 24 , p => False), (a => 40 , b => 56 , p => False), (a => 4  , b => 20 , p => False), (a => 36 , b => 52 , p => False), (a => 12 , b => 28 , p => False), (a => 44 , b => 60 , p => False), (a => 2  , b => 18 , p => False), (a => 34 , b => 50 , p => False), (a => 10 , b => 26 , p => False), (a => 42 , b => 58 , p => False), (a => 6  , b => 22 , p => False), (a => 38 , b => 54 , p => False), (a => 14 , b => 30 , p => False), (a => 46 , b => 62 , p => False), (a => 1  , b => 17 , p => False), (a => 33 , b => 49 , p => False), (a => 9  , b => 25 , p => False), (a => 41 , b => 57 , p => False), (a => 5  , b => 21 , p => False), (a => 37 , b => 53 , p => False), (a => 13 , b => 29 , p => False), (a => 45 , b => 61 , p => False), (a => 3  , b => 19 , p => False), (a => 35 , b => 51 , p => False), (a => 11 , b => 27 , p => False), (a => 43 , b => 59 , p => False), (a => 7  , b => 23 , p => False), (a => 39 , b => 55 , p => False), (a => 0  , b => 63 , p => True ), (a => 15 , b => 48 , p => True ), (a => 16 , b => 47 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 40 , b => 48 , p => False), (a => 12 , b => 20 , p => False), (a => 44 , b => 52 , p => False), (a => 10 , b => 18 , p => False), (a => 42 , b => 50 , p => False), (a => 14 , b => 22 , p => False), (a => 46 , b => 54 , p => False), (a => 9  , b => 17 , p => False), (a => 41 , b => 49 , p => False), (a => 13 , b => 21 , p => False), (a => 45 , b => 53 , p => False), (a => 11 , b => 19 , p => False), (a => 43 , b => 51 , p => False), (a => 15 , b => 23 , p => False), (a => 47 , b => 55 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 2  , b => 61 , p => True ), (a => 3  , b => 60 , p => True ), (a => 4  , b => 59 , p => True ), (a => 5  , b => 58 , p => True ), (a => 6  , b => 57 , p => True ), (a => 7  , b => 56 , p => True ), (a => 24 , b => 39 , p => True ), (a => 25 , b => 38 , p => True ), (a => 26 , b => 37 , p => True ), (a => 27 , b => 36 , p => True ), (a => 28 , b => 35 , p => True ), (a => 29 , b => 34 , p => True ), (a => 30 , b => 33 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 36 , b => 40 , p => False), (a => 44 , b => 48 , p => False), (a => 52 , b => 56 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 38 , b => 42 , p => False), (a => 46 , b => 50 , p => False), (a => 54 , b => 58 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 37 , b => 41 , p => False), (a => 45 , b => 49 , p => False), (a => 53 , b => 57 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 39 , b => 43 , p => False), (a => 47 , b => 51 , p => False), (a => 55 , b => 59 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 2  , b => 61 , p => True ), (a => 3  , b => 60 , p => True ), (a => 28 , b => 35 , p => True ), (a => 29 , b => 34 , p => True ), (a => 30 , b => 33 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 46 , b => 48 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 47 , b => 49 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 26 , b => 61 , p => True ), (a => 27 , b => 60 , p => True ), (a => 28 , b => 59 , p => True ), (a => 29 , b => 58 , p => True ), (a => 30 , b => 33 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 47 , b => 48 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 0  , b => 63 , p => True ), (a => 25 , b => 62 , p => True ), (a => 26 , b => 61 , p => True ), (a => 27 , b => 60 , p => True ), (a => 28 , b => 59 , p => True ), (a => 29 , b => 58 , p => True ), (a => 30 , b => 57 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 16 , b => 48 , p => False), (a => 8  , b => 40 , p => False), (a => 4  , b => 36 , p => False), (a => 20 , b => 52 , p => False), (a => 12 , b => 44 , p => False), (a => 2  , b => 34 , p => False), (a => 18 , b => 50 , p => False), (a => 10 , b => 42 , p => False), (a => 6  , b => 38 , p => False), (a => 22 , b => 54 , p => False), (a => 14 , b => 46 , p => False), (a => 1  , b => 33 , p => False), (a => 17 , b => 49 , p => False), (a => 9  , b => 41 , p => False), (a => 5  , b => 37 , p => False), (a => 21 , b => 53 , p => False), (a => 13 , b => 45 , p => False), (a => 3  , b => 35 , p => False), (a => 19 , b => 51 , p => False), (a => 11 , b => 43 , p => False), (a => 7  , b => 39 , p => False), (a => 23 , b => 55 , p => False), (a => 15 , b => 47 , p => False), (a => 0  , b => 63 , p => True ), (a => 24 , b => 62 , p => True ), (a => 25 , b => 61 , p => True ), (a => 26 , b => 60 , p => True ), (a => 27 , b => 59 , p => True ), (a => 28 , b => 58 , p => True ), (a => 29 , b => 57 , p => True ), (a => 30 , b => 56 , p => True ), (a => 31 , b => 32 , p => True )),
                    ((a => 16 , b => 32 , p => False), (a => 20 , b => 36 , p => False), (a => 18 , b => 34 , p => False), (a => 22 , b => 38 , p => False), (a => 17 , b => 33 , p => False), (a => 21 , b => 37 , p => False), (a => 19 , b => 35 , p => False), (a => 23 , b => 39 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 2  , b => 61 , p => True ), (a => 3  , b => 60 , p => True ), (a => 4  , b => 59 , p => True ), (a => 5  , b => 58 , p => True ), (a => 6  , b => 57 , p => True ), (a => 7  , b => 56 , p => True ), (a => 8  , b => 55 , p => True ), (a => 9  , b => 54 , p => True ), (a => 10 , b => 53 , p => True ), (a => 11 , b => 52 , p => True ), (a => 12 , b => 51 , p => True ), (a => 13 , b => 50 , p => True ), (a => 14 , b => 49 , p => True ), (a => 15 , b => 48 , p => True ), (a => 24 , b => 47 , p => True ), (a => 25 , b => 46 , p => True ), (a => 26 , b => 45 , p => True ), (a => 27 , b => 44 , p => True ), (a => 28 , b => 43 , p => True ), (a => 29 , b => 42 , p => True ), (a => 30 , b => 41 , p => True ), (a => 31 , b => 40 , p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 12 , b => 20 , p => False), (a => 10 , b => 18 , p => False), (a => 14 , b => 22 , p => False), (a => 9  , b => 17 , p => False), (a => 13 , b => 21 , p => False), (a => 11 , b => 19 , p => False), (a => 15 , b => 23 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 2  , b => 61 , p => True ), (a => 3  , b => 60 , p => True ), (a => 4  , b => 59 , p => True ), (a => 5  , b => 58 , p => True ), (a => 6  , b => 57 , p => True ), (a => 7  , b => 56 , p => True ), (a => 24 , b => 55 , p => True ), (a => 25 , b => 54 , p => True ), (a => 26 , b => 53 , p => True ), (a => 27 , b => 52 , p => True ), (a => 28 , b => 51 , p => True ), (a => 29 , b => 50 , p => True ), (a => 30 , b => 49 , p => True ), (a => 31 , b => 48 , p => True ), (a => 32 , b => 47 , p => True ), (a => 33 , b => 46 , p => True ), (a => 34 , b => 45 , p => True ), (a => 35 , b => 44 , p => True ), (a => 36 , b => 43 , p => True ), (a => 37 , b => 42 , p => True ), (a => 38 , b => 41 , p => True ), (a => 39 , b => 40 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 2  , b => 61 , p => True ), (a => 3  , b => 60 , p => True ), (a => 20 , b => 59 , p => True ), (a => 21 , b => 58 , p => True ), (a => 22 , b => 57 , p => True ), (a => 23 , b => 56 , p => True ), (a => 24 , b => 55 , p => True ), (a => 25 , b => 54 , p => True ), (a => 26 , b => 53 , p => True ), (a => 27 , b => 52 , p => True ), (a => 28 , b => 51 , p => True ), (a => 29 , b => 50 , p => True ), (a => 30 , b => 49 , p => True ), (a => 31 , b => 48 , p => True ), (a => 32 , b => 47 , p => True ), (a => 33 , b => 46 , p => True ), (a => 34 , b => 45 , p => True ), (a => 35 , b => 44 , p => True ), (a => 36 , b => 43 , p => True ), (a => 37 , b => 42 , p => True ), (a => 38 , b => 41 , p => True ), (a => 39 , b => 40 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 0  , b => 63 , p => True ), (a => 1  , b => 62 , p => True ), (a => 18 , b => 61 , p => True ), (a => 19 , b => 60 , p => True ), (a => 20 , b => 59 , p => True ), (a => 21 , b => 58 , p => True ), (a => 22 , b => 57 , p => True ), (a => 23 , b => 56 , p => True ), (a => 24 , b => 55 , p => True ), (a => 25 , b => 54 , p => True ), (a => 26 , b => 53 , p => True ), (a => 27 , b => 52 , p => True ), (a => 28 , b => 51 , p => True ), (a => 29 , b => 50 , p => True ), (a => 30 , b => 49 , p => True ), (a => 31 , b => 48 , p => True ), (a => 32 , b => 47 , p => True ), (a => 33 , b => 46 , p => True ), (a => 34 , b => 45 , p => True ), (a => 35 , b => 44 , p => True ), (a => 36 , b => 43 , p => True ), (a => 37 , b => 42 , p => True ), (a => 38 , b => 41 , p => True ), (a => 39 , b => 40 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 0  , b => 63 , p => True ), (a => 17 , b => 62 , p => True ), (a => 18 , b => 61 , p => True ), (a => 19 , b => 60 , p => True ), (a => 20 , b => 59 , p => True ), (a => 21 , b => 58 , p => True ), (a => 22 , b => 57 , p => True ), (a => 23 , b => 56 , p => True ), (a => 24 , b => 55 , p => True ), (a => 25 , b => 54 , p => True ), (a => 26 , b => 53 , p => True ), (a => 27 , b => 52 , p => True ), (a => 28 , b => 51 , p => True ), (a => 29 , b => 50 , p => True ), (a => 30 , b => 49 , p => True ), (a => 31 , b => 48 , p => True ), (a => 32 , b => 47 , p => True ), (a => 33 , b => 46 , p => True ), (a => 34 , b => 45 , p => True ), (a => 35 , b => 44 , p => True ), (a => 36 , b => 43 , p => True ), (a => 37 , b => 42 , p => True ), (a => 38 , b => 41 , p => True ), (a => 39 , b => 40 , p => True ))
                    );

            when 88 => return (
                    ((a => 0  , b => 1  , p => False), (a => 2  , b => 3  , p => False), (a => 4  , b => 5  , p => False), (a => 6  , b => 7  , p => False), (a => 8  , b => 9  , p => False), (a => 10 , b => 11 , p => False), (a => 12 , b => 13 , p => False), (a => 14 , b => 15 , p => False), (a => 16 , b => 17 , p => False), (a => 18 , b => 19 , p => False), (a => 20 , b => 21 , p => False), (a => 22 , b => 23 , p => False), (a => 24 , b => 25 , p => False), (a => 26 , b => 27 , p => False), (a => 28 , b => 29 , p => False), (a => 30 , b => 31 , p => False), (a => 32 , b => 33 , p => False), (a => 34 , b => 35 , p => False), (a => 36 , b => 37 , p => False), (a => 38 , b => 39 , p => False), (a => 40 , b => 41 , p => False), (a => 42 , b => 43 , p => False), (a => 44 , b => 45 , p => False), (a => 46 , b => 47 , p => False), (a => 48 , b => 49 , p => False), (a => 50 , b => 51 , p => False), (a => 52 , b => 53 , p => False), (a => 54 , b => 55 , p => False), (a => 56 , b => 57 , p => False), (a => 58 , b => 59 , p => False), (a => 60 , b => 61 , p => False), (a => 62 , b => 63 , p => False), (a => 64 , b => 65 , p => False), (a => 66 , b => 67 , p => False), (a => 68 , b => 69 , p => False), (a => 70 , b => 71 , p => False), (a => 72 , b => 73 , p => False), (a => 74 , b => 75 , p => False), (a => 76 , b => 77 , p => False), (a => 78 , b => 79 , p => False), (a => 80 , b => 81 , p => False), (a => 82 , b => 83 , p => False), (a => 84 , b => 85 , p => False), (a => 86 , b => 87 , p => False)),
                    ((a => 0  , b => 2  , p => False), (a => 4  , b => 6  , p => False), (a => 8  , b => 10 , p => False), (a => 12 , b => 14 , p => False), (a => 16 , b => 18 , p => False), (a => 20 , b => 22 , p => False), (a => 24 , b => 26 , p => False), (a => 28 , b => 30 , p => False), (a => 32 , b => 34 , p => False), (a => 36 , b => 38 , p => False), (a => 40 , b => 42 , p => False), (a => 44 , b => 46 , p => False), (a => 48 , b => 50 , p => False), (a => 52 , b => 54 , p => False), (a => 56 , b => 58 , p => False), (a => 60 , b => 62 , p => False), (a => 64 , b => 66 , p => False), (a => 68 , b => 70 , p => False), (a => 72 , b => 74 , p => False), (a => 76 , b => 78 , p => False), (a => 80 , b => 82 , p => False), (a => 84 , b => 86 , p => False), (a => 1  , b => 3  , p => False), (a => 5  , b => 7  , p => False), (a => 9  , b => 11 , p => False), (a => 13 , b => 15 , p => False), (a => 17 , b => 19 , p => False), (a => 21 , b => 23 , p => False), (a => 25 , b => 27 , p => False), (a => 29 , b => 31 , p => False), (a => 33 , b => 35 , p => False), (a => 37 , b => 39 , p => False), (a => 41 , b => 43 , p => False), (a => 45 , b => 47 , p => False), (a => 49 , b => 51 , p => False), (a => 53 , b => 55 , p => False), (a => 57 , b => 59 , p => False), (a => 61 , b => 63 , p => False), (a => 65 , b => 67 , p => False), (a => 69 , b => 71 , p => False), (a => 73 , b => 75 , p => False), (a => 77 , b => 79 , p => False), (a => 81 , b => 83 , p => False), (a => 85 , b => 87 , p => False)),
                    ((a => 1  , b => 2  , p => False), (a => 5  , b => 6  , p => False), (a => 9  , b => 10 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 21 , b => 22 , p => False), (a => 25 , b => 26 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 37 , b => 38 , p => False), (a => 41 , b => 42 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 53 , b => 54 , p => False), (a => 57 , b => 58 , p => False), (a => 61 , b => 62 , p => False), (a => 65 , b => 66 , p => False), (a => 69 , b => 70 , p => False), (a => 73 , b => 74 , p => False), (a => 77 , b => 78 , p => False), (a => 81 , b => 82 , p => False), (a => 85 , b => 86 , p => False), (a => 0  , b => 4  , p => False), (a => 8  , b => 12 , p => False), (a => 16 , b => 20 , p => False), (a => 24 , b => 28 , p => False), (a => 32 , b => 36 , p => False), (a => 40 , b => 44 , p => False), (a => 48 , b => 52 , p => False), (a => 56 , b => 60 , p => False), (a => 64 , b => 68 , p => False), (a => 72 , b => 76 , p => False), (a => 80 , b => 84 , p => False), (a => 3  , b => 7  , p => False), (a => 11 , b => 15 , p => False), (a => 19 , b => 23 , p => False), (a => 27 , b => 31 , p => False), (a => 35 , b => 39 , p => False), (a => 43 , b => 47 , p => False), (a => 51 , b => 55 , p => False), (a => 59 , b => 63 , p => False), (a => 67 , b => 71 , p => False), (a => 75 , b => 79 , p => False), (a => 83 , b => 87 , p => False)),
                    ((a => 2  , b => 6  , p => False), (a => 10 , b => 14 , p => False), (a => 18 , b => 22 , p => False), (a => 26 , b => 30 , p => False), (a => 34 , b => 38 , p => False), (a => 42 , b => 46 , p => False), (a => 50 , b => 54 , p => False), (a => 58 , b => 62 , p => False), (a => 66 , b => 70 , p => False), (a => 74 , b => 78 , p => False), (a => 82 , b => 86 , p => False), (a => 1  , b => 5  , p => False), (a => 9  , b => 13 , p => False), (a => 17 , b => 21 , p => False), (a => 25 , b => 29 , p => False), (a => 33 , b => 37 , p => False), (a => 41 , b => 45 , p => False), (a => 49 , b => 53 , p => False), (a => 57 , b => 61 , p => False), (a => 65 , b => 69 , p => False), (a => 73 , b => 77 , p => False), (a => 81 , b => 85 , p => False), (a => 0  , b => 8  , p => False), (a => 16 , b => 24 , p => False), (a => 32 , b => 40 , p => False), (a => 48 , b => 56 , p => False), (a => 64 , b => 72 , p => False), (a => 7  , b => 15 , p => False), (a => 23 , b => 31 , p => False), (a => 39 , b => 47 , p => False), (a => 55 , b => 63 , p => False), (a => 71 , b => 79 , p => False), (a => 3  , b => 87 , p => True ), (a => 4  , b => 84 , p => True ), (a => 11 , b => 83 , p => True ), (a => 12 , b => 80 , p => True ), (a => 19 , b => 76 , p => True ), (a => 20 , b => 75 , p => True ), (a => 27 , b => 68 , p => True ), (a => 28 , b => 67 , p => True ), (a => 35 , b => 60 , p => True ), (a => 36 , b => 59 , p => True ), (a => 43 , b => 52 , p => True ), (a => 44 , b => 51 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 10 , b => 12 , p => False), (a => 18 , b => 20 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 42 , b => 44 , p => False), (a => 50 , b => 52 , p => False), (a => 58 , b => 60 , p => False), (a => 66 , b => 68 , p => False), (a => 74 , b => 76 , p => False), (a => 82 , b => 84 , p => False), (a => 3  , b => 5  , p => False), (a => 11 , b => 13 , p => False), (a => 19 , b => 21 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 43 , b => 45 , p => False), (a => 51 , b => 53 , p => False), (a => 59 , b => 61 , p => False), (a => 67 , b => 69 , p => False), (a => 75 , b => 77 , p => False), (a => 83 , b => 85 , p => False), (a => 0  , b => 16 , p => False), (a => 32 , b => 48 , p => False), (a => 64 , b => 80 , p => False), (a => 15 , b => 31 , p => False), (a => 47 , b => 63 , p => False), (a => 1  , b => 87 , p => True ), (a => 6  , b => 86 , p => True ), (a => 7  , b => 81 , p => True ), (a => 8  , b => 79 , p => True ), (a => 9  , b => 78 , p => True ), (a => 14 , b => 73 , p => True ), (a => 17 , b => 72 , p => True ), (a => 22 , b => 71 , p => True ), (a => 23 , b => 70 , p => True ), (a => 24 , b => 65 , p => True ), (a => 25 , b => 62 , p => True ), (a => 30 , b => 57 , p => True ), (a => 33 , b => 56 , p => True ), (a => 38 , b => 55 , p => True ), (a => 39 , b => 54 , p => True ), (a => 40 , b => 49 , p => True ), (a => 41 , b => 46 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 0  , b => 32 , p => False), (a => 31 , b => 63 , p => False), (a => 7  , b => 87 , p => True ), (a => 8  , b => 80 , p => True ), (a => 15 , b => 79 , p => True ), (a => 16 , b => 72 , p => True ), (a => 23 , b => 71 , p => True ), (a => 24 , b => 64 , p => True ), (a => 39 , b => 56 , p => True ), (a => 40 , b => 55 , p => True ), (a => 47 , b => 48 , p => True )),
                    ((a => 4  , b => 12 , p => False), (a => 20 , b => 28 , p => False), (a => 36 , b => 44 , p => False), (a => 52 , b => 60 , p => False), (a => 68 , b => 76 , p => False), (a => 2  , b => 10 , p => False), (a => 18 , b => 26 , p => False), (a => 34 , b => 42 , p => False), (a => 50 , b => 58 , p => False), (a => 66 , b => 74 , p => False), (a => 6  , b => 14 , p => False), (a => 22 , b => 30 , p => False), (a => 38 , b => 46 , p => False), (a => 54 , b => 62 , p => False), (a => 70 , b => 78 , p => False), (a => 1  , b => 9  , p => False), (a => 17 , b => 25 , p => False), (a => 33 , b => 41 , p => False), (a => 49 , b => 57 , p => False), (a => 65 , b => 73 , p => False), (a => 5  , b => 13 , p => False), (a => 21 , b => 29 , p => False), (a => 37 , b => 45 , p => False), (a => 53 , b => 61 , p => False), (a => 69 , b => 77 , p => False), (a => 3  , b => 11 , p => False), (a => 19 , b => 27 , p => False), (a => 35 , b => 43 , p => False), (a => 51 , b => 59 , p => False), (a => 67 , b => 75 , p => False), (a => 0  , b => 64 , p => False), (a => 82 , b => 84 , p => False), (a => 83 , b => 85 , p => False), (a => 7  , b => 87 , p => True ), (a => 8  , b => 86 , p => True ), (a => 15 , b => 81 , p => True ), (a => 16 , b => 80 , p => True ), (a => 23 , b => 79 , p => True ), (a => 24 , b => 72 , p => True ), (a => 31 , b => 71 , p => True ), (a => 32 , b => 63 , p => True ), (a => 39 , b => 56 , p => True ), (a => 40 , b => 55 , p => True ), (a => 47 , b => 48 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 20 , b => 24 , p => False), (a => 36 , b => 40 , p => False), (a => 52 , b => 56 , p => False), (a => 68 , b => 72 , p => False), (a => 6  , b => 10 , p => False), (a => 22 , b => 26 , p => False), (a => 38 , b => 42 , p => False), (a => 54 , b => 58 , p => False), (a => 70 , b => 74 , p => False), (a => 5  , b => 9  , p => False), (a => 21 , b => 25 , p => False), (a => 37 , b => 41 , p => False), (a => 53 , b => 57 , p => False), (a => 69 , b => 73 , p => False), (a => 7  , b => 11 , p => False), (a => 23 , b => 27 , p => False), (a => 39 , b => 43 , p => False), (a => 55 , b => 59 , p => False), (a => 71 , b => 75 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 80 , p => True ), (a => 2  , b => 79 , p => True ), (a => 3  , b => 78 , p => True ), (a => 12 , b => 77 , p => True ), (a => 13 , b => 76 , p => True ), (a => 14 , b => 67 , p => True ), (a => 15 , b => 66 , p => True ), (a => 16 , b => 65 , p => True ), (a => 17 , b => 64 , p => True ), (a => 18 , b => 63 , p => True ), (a => 19 , b => 62 , p => True ), (a => 28 , b => 61 , p => True ), (a => 29 , b => 60 , p => True ), (a => 30 , b => 51 , p => True ), (a => 31 , b => 50 , p => True ), (a => 32 , b => 49 , p => True ), (a => 33 , b => 48 , p => True ), (a => 34 , b => 47 , p => True ), (a => 35 , b => 46 , p => True ), (a => 44 , b => 45 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 14 , b => 85 , p => True ), (a => 15 , b => 84 , p => True ), (a => 16 , b => 83 , p => True ), (a => 17 , b => 82 , p => True ), (a => 30 , b => 81 , p => True ), (a => 31 , b => 80 , p => True ), (a => 32 , b => 79 , p => True ), (a => 33 , b => 78 , p => True ), (a => 46 , b => 65 , p => True ), (a => 47 , b => 64 , p => True ), (a => 48 , b => 63 , p => True ), (a => 49 , b => 62 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 0  , b => 87 , p => True ), (a => 15 , b => 86 , p => True ), (a => 16 , b => 85 , p => True ), (a => 31 , b => 84 , p => True ), (a => 32 , b => 83 , p => True ), (a => 47 , b => 82 , p => True ), (a => 48 , b => 81 , p => True ), (a => 63 , b => 80 , p => True ), (a => 64 , b => 79 , p => True )),
                    ((a => 8  , b => 24 , p => False), (a => 40 , b => 56 , p => False), (a => 4  , b => 20 , p => False), (a => 36 , b => 52 , p => False), (a => 68 , b => 84 , p => False), (a => 12 , b => 28 , p => False), (a => 44 , b => 60 , p => False), (a => 2  , b => 18 , p => False), (a => 34 , b => 50 , p => False), (a => 66 , b => 82 , p => False), (a => 10 , b => 26 , p => False), (a => 42 , b => 58 , p => False), (a => 6  , b => 22 , p => False), (a => 38 , b => 54 , p => False), (a => 70 , b => 86 , p => False), (a => 14 , b => 30 , p => False), (a => 46 , b => 62 , p => False), (a => 1  , b => 17 , p => False), (a => 33 , b => 49 , p => False), (a => 65 , b => 81 , p => False), (a => 9  , b => 25 , p => False), (a => 41 , b => 57 , p => False), (a => 5  , b => 21 , p => False), (a => 37 , b => 53 , p => False), (a => 69 , b => 85 , p => False), (a => 13 , b => 29 , p => False), (a => 45 , b => 61 , p => False), (a => 3  , b => 19 , p => False), (a => 35 , b => 51 , p => False), (a => 67 , b => 83 , p => False), (a => 11 , b => 27 , p => False), (a => 43 , b => 59 , p => False), (a => 7  , b => 23 , p => False), (a => 39 , b => 55 , p => False), (a => 71 , b => 87 , p => False), (a => 72 , b => 80 , p => False), (a => 0  , b => 79 , p => True ), (a => 15 , b => 78 , p => True ), (a => 16 , b => 77 , p => True ), (a => 31 , b => 76 , p => True ), (a => 32 , b => 75 , p => True ), (a => 47 , b => 74 , p => True ), (a => 48 , b => 73 , p => True ), (a => 63 , b => 64 , p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 40 , b => 48 , p => False), (a => 12 , b => 20 , p => False), (a => 44 , b => 52 , p => False), (a => 76 , b => 84 , p => False), (a => 10 , b => 18 , p => False), (a => 42 , b => 50 , p => False), (a => 74 , b => 82 , p => False), (a => 14 , b => 22 , p => False), (a => 46 , b => 54 , p => False), (a => 78 , b => 86 , p => False), (a => 9  , b => 17 , p => False), (a => 41 , b => 49 , p => False), (a => 73 , b => 81 , p => False), (a => 13 , b => 21 , p => False), (a => 45 , b => 53 , p => False), (a => 77 , b => 85 , p => False), (a => 11 , b => 19 , p => False), (a => 43 , b => 51 , p => False), (a => 75 , b => 83 , p => False), (a => 15 , b => 23 , p => False), (a => 47 , b => 55 , p => False), (a => 79 , b => 87 , p => False), (a => 68 , b => 72 , p => False), (a => 0  , b => 80 , p => True ), (a => 1  , b => 71 , p => True ), (a => 2  , b => 70 , p => True ), (a => 3  , b => 69 , p => True ), (a => 4  , b => 67 , p => True ), (a => 5  , b => 66 , p => True ), (a => 6  , b => 65 , p => True ), (a => 7  , b => 64 , p => True ), (a => 24 , b => 63 , p => True ), (a => 25 , b => 62 , p => True ), (a => 26 , b => 61 , p => True ), (a => 27 , b => 60 , p => True ), (a => 28 , b => 59 , p => True ), (a => 29 , b => 58 , p => True ), (a => 30 , b => 57 , p => True ), (a => 31 , b => 56 , p => True ), (a => 32 , b => 39 , p => True ), (a => 33 , b => 38 , p => True ), (a => 34 , b => 37 , p => True ), (a => 35 , b => 36 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 36 , b => 40 , p => False), (a => 44 , b => 48 , p => False), (a => 52 , b => 56 , p => False), (a => 76 , b => 80 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 38 , b => 42 , p => False), (a => 46 , b => 50 , p => False), (a => 54 , b => 58 , p => False), (a => 70 , b => 74 , p => False), (a => 78 , b => 82 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 37 , b => 41 , p => False), (a => 45 , b => 49 , p => False), (a => 53 , b => 57 , p => False), (a => 69 , b => 73 , p => False), (a => 77 , b => 81 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 39 , b => 43 , p => False), (a => 47 , b => 51 , p => False), (a => 55 , b => 59 , p => False), (a => 71 , b => 75 , p => False), (a => 79 , b => 83 , p => False), (a => 66 , b => 68 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 85 , p => True ), (a => 3  , b => 84 , p => True ), (a => 28 , b => 72 , p => True ), (a => 29 , b => 67 , p => True ), (a => 30 , b => 65 , p => True ), (a => 31 , b => 64 , p => True ), (a => 32 , b => 63 , p => True ), (a => 33 , b => 62 , p => True ), (a => 34 , b => 61 , p => True ), (a => 35 , b => 60 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 46 , b => 48 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 78 , b => 80 , p => False), (a => 82 , b => 84 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 47 , b => 49 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 79 , b => 81 , p => False), (a => 83 , b => 85 , p => False), (a => 65 , b => 66 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 30 , b => 68 , p => True ), (a => 31 , b => 64 , p => True ), (a => 32 , b => 63 , p => True ), (a => 33 , b => 62 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 47 , b => 48 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 79 , b => 80 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 0  , b => 87 , p => True ), (a => 31 , b => 66 , p => True ), (a => 32 , b => 65 , p => True ), (a => 63 , b => 64 , p => True )),
                    ((a => 16 , b => 48 , p => False), (a => 8  , b => 40 , p => False), (a => 24 , b => 56 , p => False), (a => 4  , b => 36 , p => False), (a => 20 , b => 52 , p => False), (a => 12 , b => 44 , p => False), (a => 28 , b => 60 , p => False), (a => 2  , b => 34 , p => False), (a => 18 , b => 50 , p => False), (a => 10 , b => 42 , p => False), (a => 26 , b => 58 , p => False), (a => 6  , b => 38 , p => False), (a => 22 , b => 54 , p => False), (a => 14 , b => 46 , p => False), (a => 30 , b => 62 , p => False), (a => 1  , b => 33 , p => False), (a => 17 , b => 49 , p => False), (a => 9  , b => 41 , p => False), (a => 25 , b => 57 , p => False), (a => 5  , b => 37 , p => False), (a => 21 , b => 53 , p => False), (a => 13 , b => 45 , p => False), (a => 29 , b => 61 , p => False), (a => 3  , b => 35 , p => False), (a => 19 , b => 51 , p => False), (a => 11 , b => 43 , p => False), (a => 27 , b => 59 , p => False), (a => 7  , b => 39 , p => False), (a => 23 , b => 55 , p => False), (a => 15 , b => 47 , p => False), (a => 72 , b => 80 , p => False), (a => 76 , b => 84 , p => False), (a => 74 , b => 82 , p => False), (a => 78 , b => 86 , p => False), (a => 73 , b => 81 , p => False), (a => 77 , b => 85 , p => False), (a => 75 , b => 83 , p => False), (a => 79 , b => 87 , p => False), (a => 0  , b => 71 , p => True ), (a => 31 , b => 70 , p => True ), (a => 32 , b => 69 , p => True ), (a => 63 , b => 68 , p => True ), (a => 64 , b => 67 , p => True ), (a => 65 , b => 66 , p => True )),
                    ((a => 16 , b => 32 , p => False), (a => 24 , b => 40 , p => False), (a => 20 , b => 36 , p => False), (a => 28 , b => 44 , p => False), (a => 18 , b => 34 , p => False), (a => 26 , b => 42 , p => False), (a => 22 , b => 38 , p => False), (a => 30 , b => 46 , p => False), (a => 17 , b => 33 , p => False), (a => 25 , b => 41 , p => False), (a => 21 , b => 37 , p => False), (a => 29 , b => 45 , p => False), (a => 19 , b => 35 , p => False), (a => 27 , b => 43 , p => False), (a => 23 , b => 39 , p => False), (a => 31 , b => 47 , p => False), (a => 68 , b => 72 , p => False), (a => 76 , b => 80 , p => False), (a => 70 , b => 74 , p => False), (a => 78 , b => 82 , p => False), (a => 69 , b => 73 , p => False), (a => 77 , b => 81 , p => False), (a => 71 , b => 75 , p => False), (a => 79 , b => 83 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 85 , p => True ), (a => 3  , b => 84 , p => True ), (a => 4  , b => 67 , p => True ), (a => 5  , b => 66 , p => True ), (a => 6  , b => 65 , p => True ), (a => 7  , b => 64 , p => True ), (a => 8  , b => 63 , p => True ), (a => 9  , b => 62 , p => True ), (a => 10 , b => 61 , p => True ), (a => 11 , b => 60 , p => True ), (a => 12 , b => 59 , p => True ), (a => 13 , b => 58 , p => True ), (a => 14 , b => 57 , p => True ), (a => 15 , b => 56 , p => True ), (a => 48 , b => 55 , p => True ), (a => 49 , b => 54 , p => True ), (a => 50 , b => 53 , p => True ), (a => 51 , b => 52 , p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 24 , b => 32 , p => False), (a => 40 , b => 48 , p => False), (a => 12 , b => 20 , p => False), (a => 28 , b => 36 , p => False), (a => 10 , b => 18 , p => False), (a => 26 , b => 34 , p => False), (a => 42 , b => 50 , p => False), (a => 14 , b => 22 , p => False), (a => 30 , b => 38 , p => False), (a => 9  , b => 17 , p => False), (a => 25 , b => 33 , p => False), (a => 41 , b => 49 , p => False), (a => 13 , b => 21 , p => False), (a => 29 , b => 37 , p => False), (a => 11 , b => 19 , p => False), (a => 27 , b => 35 , p => False), (a => 43 , b => 51 , p => False), (a => 15 , b => 23 , p => False), (a => 31 , b => 39 , p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 78 , b => 80 , p => False), (a => 82 , b => 84 , p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 79 , b => 81 , p => False), (a => 83 , b => 85 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 65 , p => True ), (a => 3  , b => 64 , p => True ), (a => 4  , b => 63 , p => True ), (a => 5  , b => 62 , p => True ), (a => 6  , b => 61 , p => True ), (a => 7  , b => 60 , p => True ), (a => 44 , b => 59 , p => True ), (a => 45 , b => 58 , p => True ), (a => 46 , b => 57 , p => True ), (a => 47 , b => 56 , p => True ), (a => 52 , b => 55 , p => True ), (a => 53 , b => 54 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 28 , b => 32 , p => False), (a => 36 , b => 40 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 30 , b => 34 , p => False), (a => 38 , b => 42 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 29 , b => 33 , p => False), (a => 37 , b => 41 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 31 , b => 35 , p => False), (a => 39 , b => 43 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 79 , b => 80 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 64 , p => True ), (a => 2  , b => 63 , p => True ), (a => 3  , b => 62 , p => True ), (a => 44 , b => 61 , p => True ), (a => 45 , b => 60 , p => True ), (a => 46 , b => 59 , p => True ), (a => 47 , b => 58 , p => True ), (a => 48 , b => 57 , p => True ), (a => 49 , b => 56 , p => True ), (a => 50 , b => 55 , p => True ), (a => 51 , b => 54 , p => True ), (a => 52 , b => 53 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 30 , b => 32 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 31 , b => 33 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 26 , b => 85 , p => True ), (a => 27 , b => 84 , p => True ), (a => 28 , b => 83 , p => True ), (a => 29 , b => 82 , p => True ), (a => 42 , b => 81 , p => True ), (a => 43 , b => 80 , p => True ), (a => 44 , b => 79 , p => True ), (a => 45 , b => 78 , p => True ), (a => 46 , b => 77 , p => True ), (a => 47 , b => 76 , p => True ), (a => 48 , b => 75 , p => True ), (a => 49 , b => 74 , p => True ), (a => 50 , b => 73 , p => True ), (a => 51 , b => 72 , p => True ), (a => 52 , b => 71 , p => True ), (a => 53 , b => 70 , p => True ), (a => 54 , b => 69 , p => True ), (a => 55 , b => 68 , p => True ), (a => 56 , b => 67 , p => True ), (a => 57 , b => 66 , p => True ), (a => 58 , b => 65 , p => True ), (a => 59 , b => 64 , p => True ), (a => 60 , b => 63 , p => True ), (a => 61 , b => 62 , p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 31 , b => 32 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 0  , b => 87 , p => True ), (a => 25 , b => 86 , p => True ), (a => 26 , b => 85 , p => True ), (a => 27 , b => 84 , p => True ), (a => 28 , b => 83 , p => True ), (a => 29 , b => 82 , p => True ), (a => 30 , b => 81 , p => True ), (a => 41 , b => 80 , p => True ), (a => 42 , b => 79 , p => True ), (a => 43 , b => 78 , p => True ), (a => 44 , b => 77 , p => True ), (a => 45 , b => 76 , p => True ), (a => 46 , b => 75 , p => True ), (a => 47 , b => 74 , p => True ), (a => 48 , b => 73 , p => True ), (a => 49 , b => 72 , p => True ), (a => 50 , b => 71 , p => True ), (a => 51 , b => 70 , p => True ), (a => 52 , b => 69 , p => True ), (a => 53 , b => 68 , p => True ), (a => 54 , b => 67 , p => True ), (a => 55 , b => 66 , p => True ), (a => 56 , b => 65 , p => True ), (a => 57 , b => 64 , p => True ), (a => 58 , b => 63 , p => True ), (a => 59 , b => 62 , p => True ), (a => 60 , b => 61 , p => True )),
                    ((a => 16 , b => 80 , p => False), (a => 8  , b => 72 , p => False), (a => 4  , b => 68 , p => False), (a => 20 , b => 84 , p => False), (a => 12 , b => 76 , p => False), (a => 2  , b => 66 , p => False), (a => 18 , b => 82 , p => False), (a => 10 , b => 74 , p => False), (a => 6  , b => 70 , p => False), (a => 22 , b => 86 , p => False), (a => 14 , b => 78 , p => False), (a => 1  , b => 65 , p => False), (a => 17 , b => 81 , p => False), (a => 9  , b => 73 , p => False), (a => 5  , b => 69 , p => False), (a => 21 , b => 85 , p => False), (a => 13 , b => 77 , p => False), (a => 3  , b => 67 , p => False), (a => 19 , b => 83 , p => False), (a => 11 , b => 75 , p => False), (a => 7  , b => 71 , p => False), (a => 23 , b => 87 , p => False), (a => 15 , b => 79 , p => False), (a => 32 , b => 64 , p => False), (a => 0  , b => 63 , p => True ), (a => 24 , b => 62 , p => True ), (a => 25 , b => 61 , p => True ), (a => 26 , b => 60 , p => True ), (a => 27 , b => 59 , p => True ), (a => 28 , b => 58 , p => True ), (a => 29 , b => 57 , p => True ), (a => 30 , b => 56 , p => True ), (a => 31 , b => 55 , p => True ), (a => 33 , b => 54 , p => True ), (a => 34 , b => 53 , p => True ), (a => 35 , b => 52 , p => True ), (a => 36 , b => 51 , p => True ), (a => 37 , b => 50 , p => True ), (a => 38 , b => 49 , p => True ), (a => 39 , b => 48 , p => True ), (a => 40 , b => 47 , p => True ), (a => 41 , b => 46 , p => True ), (a => 42 , b => 45 , p => True ), (a => 43 , b => 44 , p => True )),
                    ((a => 36 , b => 68 , p => False), (a => 34 , b => 66 , p => False), (a => 38 , b => 70 , p => False), (a => 33 , b => 65 , p => False), (a => 37 , b => 69 , p => False), (a => 35 , b => 67 , p => False), (a => 39 , b => 71 , p => False), (a => 16 , b => 32 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 85 , p => True ), (a => 3  , b => 84 , p => True ), (a => 4  , b => 83 , p => True ), (a => 5  , b => 82 , p => True ), (a => 6  , b => 81 , p => True ), (a => 7  , b => 80 , p => True ), (a => 8  , b => 79 , p => True ), (a => 9  , b => 78 , p => True ), (a => 10 , b => 77 , p => True ), (a => 11 , b => 76 , p => True ), (a => 12 , b => 75 , p => True ), (a => 13 , b => 74 , p => True ), (a => 14 , b => 73 , p => True ), (a => 15 , b => 72 , p => True ), (a => 17 , b => 64 , p => True ), (a => 18 , b => 63 , p => True ), (a => 19 , b => 62 , p => True ), (a => 20 , b => 61 , p => True ), (a => 21 , b => 60 , p => True ), (a => 22 , b => 59 , p => True ), (a => 23 , b => 58 , p => True ), (a => 24 , b => 57 , p => True ), (a => 25 , b => 56 , p => True ), (a => 26 , b => 55 , p => True ), (a => 27 , b => 54 , p => True ), (a => 28 , b => 53 , p => True ), (a => 29 , b => 52 , p => True ), (a => 30 , b => 51 , p => True ), (a => 31 , b => 50 , p => True ), (a => 40 , b => 49 , p => True ), (a => 41 , b => 48 , p => True ), (a => 42 , b => 47 , p => True ), (a => 43 , b => 46 , p => True ), (a => 44 , b => 45 , p => True )),
                    ((a => 20 , b => 36 , p => False), (a => 18 , b => 34 , p => False), (a => 22 , b => 38 , p => False), (a => 17 , b => 33 , p => False), (a => 21 , b => 37 , p => False), (a => 19 , b => 35 , p => False), (a => 23 , b => 39 , p => False), (a => 8  , b => 16 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 85 , p => True ), (a => 3  , b => 84 , p => True ), (a => 4  , b => 83 , p => True ), (a => 5  , b => 82 , p => True ), (a => 6  , b => 81 , p => True ), (a => 7  , b => 80 , p => True ), (a => 9  , b => 79 , p => True ), (a => 10 , b => 78 , p => True ), (a => 11 , b => 77 , p => True ), (a => 12 , b => 76 , p => True ), (a => 13 , b => 75 , p => True ), (a => 14 , b => 74 , p => True ), (a => 15 , b => 73 , p => True ), (a => 24 , b => 72 , p => True ), (a => 25 , b => 71 , p => True ), (a => 26 , b => 70 , p => True ), (a => 27 , b => 69 , p => True ), (a => 28 , b => 68 , p => True ), (a => 29 , b => 67 , p => True ), (a => 30 , b => 66 , p => True ), (a => 31 , b => 65 , p => True ), (a => 32 , b => 64 , p => True ), (a => 40 , b => 63 , p => True ), (a => 41 , b => 62 , p => True ), (a => 42 , b => 61 , p => True ), (a => 43 , b => 60 , p => True ), (a => 44 , b => 59 , p => True ), (a => 45 , b => 58 , p => True ), (a => 46 , b => 57 , p => True ), (a => 47 , b => 56 , p => True ), (a => 48 , b => 55 , p => True ), (a => 49 , b => 54 , p => True ), (a => 50 , b => 53 , p => True ), (a => 51 , b => 52 , p => True )),
                    ((a => 12 , b => 20 , p => False), (a => 10 , b => 18 , p => False), (a => 14 , b => 22 , p => False), (a => 9  , b => 17 , p => False), (a => 13 , b => 21 , p => False), (a => 11 , b => 19 , p => False), (a => 15 , b => 23 , p => False), (a => 4  , b => 8  , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 85 , p => True ), (a => 3  , b => 84 , p => True ), (a => 5  , b => 83 , p => True ), (a => 6  , b => 82 , p => True ), (a => 7  , b => 81 , p => True ), (a => 16 , b => 80 , p => True ), (a => 24 , b => 79 , p => True ), (a => 25 , b => 78 , p => True ), (a => 26 , b => 77 , p => True ), (a => 27 , b => 76 , p => True ), (a => 28 , b => 75 , p => True ), (a => 29 , b => 74 , p => True ), (a => 30 , b => 73 , p => True ), (a => 31 , b => 72 , p => True ), (a => 32 , b => 71 , p => True ), (a => 33 , b => 70 , p => True ), (a => 34 , b => 69 , p => True ), (a => 35 , b => 68 , p => True ), (a => 36 , b => 67 , p => True ), (a => 37 , b => 66 , p => True ), (a => 38 , b => 65 , p => True ), (a => 39 , b => 64 , p => True ), (a => 40 , b => 63 , p => True ), (a => 41 , b => 62 , p => True ), (a => 42 , b => 61 , p => True ), (a => 43 , b => 60 , p => True ), (a => 44 , b => 59 , p => True ), (a => 45 , b => 58 , p => True ), (a => 46 , b => 57 , p => True ), (a => 47 , b => 56 , p => True ), (a => 48 , b => 55 , p => True ), (a => 49 , b => 54 , p => True ), (a => 50 , b => 53 , p => True ), (a => 51 , b => 52 , p => True )),
                    ((a => 12 , b => 16 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 2  , b => 4  , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 3  , b => 85 , p => True ), (a => 8  , b => 84 , p => True ), (a => 20 , b => 83 , p => True ), (a => 21 , b => 82 , p => True ), (a => 22 , b => 81 , p => True ), (a => 23 , b => 80 , p => True ), (a => 24 , b => 79 , p => True ), (a => 25 , b => 78 , p => True ), (a => 26 , b => 77 , p => True ), (a => 27 , b => 76 , p => True ), (a => 28 , b => 75 , p => True ), (a => 29 , b => 74 , p => True ), (a => 30 , b => 73 , p => True ), (a => 31 , b => 72 , p => True ), (a => 32 , b => 71 , p => True ), (a => 33 , b => 70 , p => True ), (a => 34 , b => 69 , p => True ), (a => 35 , b => 68 , p => True ), (a => 36 , b => 67 , p => True ), (a => 37 , b => 66 , p => True ), (a => 38 , b => 65 , p => True ), (a => 39 , b => 64 , p => True ), (a => 40 , b => 63 , p => True ), (a => 41 , b => 62 , p => True ), (a => 42 , b => 61 , p => True ), (a => 43 , b => 60 , p => True ), (a => 44 , b => 59 , p => True ), (a => 45 , b => 58 , p => True ), (a => 46 , b => 57 , p => True ), (a => 47 , b => 56 , p => True ), (a => 48 , b => 55 , p => True ), (a => 49 , b => 54 , p => True ), (a => 50 , b => 53 , p => True ), (a => 51 , b => 52 , p => True )),
                    ((a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 1  , b => 2  , p => False), (a => 0  , b => 87 , p => True ), (a => 4  , b => 86 , p => True ), (a => 18 , b => 85 , p => True ), (a => 19 , b => 84 , p => True ), (a => 20 , b => 83 , p => True ), (a => 21 , b => 82 , p => True ), (a => 22 , b => 81 , p => True ), (a => 23 , b => 80 , p => True ), (a => 24 , b => 79 , p => True ), (a => 25 , b => 78 , p => True ), (a => 26 , b => 77 , p => True ), (a => 27 , b => 76 , p => True ), (a => 28 , b => 75 , p => True ), (a => 29 , b => 74 , p => True ), (a => 30 , b => 73 , p => True ), (a => 31 , b => 72 , p => True ), (a => 32 , b => 71 , p => True ), (a => 33 , b => 70 , p => True ), (a => 34 , b => 69 , p => True ), (a => 35 , b => 68 , p => True ), (a => 36 , b => 67 , p => True ), (a => 37 , b => 66 , p => True ), (a => 38 , b => 65 , p => True ), (a => 39 , b => 64 , p => True ), (a => 40 , b => 63 , p => True ), (a => 41 , b => 62 , p => True ), (a => 42 , b => 61 , p => True ), (a => 43 , b => 60 , p => True ), (a => 44 , b => 59 , p => True ), (a => 45 , b => 58 , p => True ), (a => 46 , b => 57 , p => True ), (a => 47 , b => 56 , p => True ), (a => 48 , b => 55 , p => True ), (a => 49 , b => 54 , p => True ), (a => 50 , b => 53 , p => True ), (a => 51 , b => 52 , p => True )),
                    ((a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 0  , b => 87 , p => True ), (a => 1  , b => 86 , p => True ), (a => 2  , b => 85 , p => True ), (a => 17 , b => 84 , p => True ), (a => 18 , b => 83 , p => True ), (a => 19 , b => 82 , p => True ), (a => 20 , b => 81 , p => True ), (a => 21 , b => 80 , p => True ), (a => 22 , b => 79 , p => True ), (a => 23 , b => 78 , p => True ), (a => 24 , b => 77 , p => True ), (a => 25 , b => 76 , p => True ), (a => 26 , b => 75 , p => True ), (a => 27 , b => 74 , p => True ), (a => 28 , b => 73 , p => True ), (a => 29 , b => 72 , p => True ), (a => 30 , b => 71 , p => True ), (a => 31 , b => 70 , p => True ), (a => 32 , b => 69 , p => True ), (a => 33 , b => 68 , p => True ), (a => 34 , b => 67 , p => True ), (a => 35 , b => 66 , p => True ), (a => 36 , b => 65 , p => True ), (a => 37 , b => 64 , p => True ), (a => 38 , b => 63 , p => True ), (a => 39 , b => 62 , p => True ), (a => 40 , b => 61 , p => True ), (a => 41 , b => 60 , p => True ), (a => 42 , b => 59 , p => True ), (a => 43 , b => 58 , p => True ), (a => 44 , b => 57 , p => True ), (a => 45 , b => 56 , p => True ), (a => 46 , b => 55 , p => True ), (a => 47 , b => 54 , p => True ), (a => 48 , b => 53 , p => True ), (a => 49 , b => 52 , p => True ), (a => 50 , b => 51 , p => True ))
                    );

					
			
			when 352 => return (
                    ((a => 0  , b => 2  , p => False), (a => 4  , b => 6  , p => False), (a => 8  , b => 10 , p => False), (a => 12 , b => 14 , p => False), (a => 16 , b => 18 , p => False), (a => 20 , b => 22 , p => False), (a => 24 , b => 26 , p => False), (a => 28 , b => 30 , p => False), (a => 32 , b => 34 , p => False), (a => 36 , b => 38 , p => False), (a => 40 , b => 42 , p => False), (a => 44 , b => 46 , p => False), (a => 48 , b => 50 , p => False), (a => 52 , b => 54 , p => False), (a => 56 , b => 58 , p => False), (a => 60 , b => 62 , p => False), (a => 1  , b => 3  , p => False), (a => 5  , b => 7  , p => False), (a => 9  , b => 11 , p => False), (a => 13 , b => 15 , p => False), (a => 17 , b => 19 , p => False), (a => 21 , b => 23 , p => False), (a => 25 , b => 27 , p => False), (a => 29 , b => 31 , p => False), (a => 33 , b => 35 , p => False), (a => 37 , b => 39 , p => False), (a => 41 , b => 43 , p => False), (a => 45 , b => 47 , p => False), (a => 49 , b => 51 , p => False), (a => 53 , b => 55 , p => False), (a => 57 , b => 59 , p => False), (a => 61 , b => 63 , p => False), (a => 64 , b => 68 , p => False), (a => 72 , b => 76 , p => False), (a => 80 , b => 84 , p => False), (a => 88 , b => 92 , p => False), (a => 96 , b => 100, p => False), (a => 104, b => 108, p => False), (a => 112, b => 116, p => False), (a => 120, b => 124, p => False), (a => 128, b => 132, p => False), (a => 136, b => 140, p => False), (a => 144, b => 148, p => False), (a => 152, b => 156, p => False), (a => 160, b => 164, p => False), (a => 168, b => 172, p => False), (a => 176, b => 180, p => False), (a => 184, b => 188, p => False), (a => 192, b => 196, p => False), (a => 200, b => 204, p => False), (a => 208, b => 212, p => False), (a => 216, b => 220, p => False), (a => 224, b => 228, p => False), (a => 232, b => 236, p => False), (a => 240, b => 244, p => False), (a => 248, b => 252, p => False), (a => 256, b => 260, p => False), (a => 264, b => 268, p => False), (a => 272, b => 276, p => False), (a => 280, b => 284, p => False), (a => 288, b => 292, p => False), (a => 296, b => 300, p => False), (a => 304, b => 308, p => False), (a => 312, b => 316, p => False), (a => 320, b => 324, p => False), (a => 328, b => 332, p => False), (a => 336, b => 340, p => False), (a => 344, b => 348, p => False), (a => 67 , b => 71 , p => False), (a => 75 , b => 79 , p => False), (a => 83 , b => 87 , p => False), (a => 91 , b => 95 , p => False), (a => 99 , b => 103, p => False), (a => 107, b => 111, p => False), (a => 115, b => 119, p => False), (a => 123, b => 127, p => False), (a => 131, b => 135, p => False), (a => 139, b => 143, p => False), (a => 147, b => 151, p => False), (a => 155, b => 159, p => False), (a => 163, b => 167, p => False), (a => 171, b => 175, p => False), (a => 179, b => 183, p => False), (a => 187, b => 191, p => False), (a => 195, b => 199, p => False), (a => 203, b => 207, p => False), (a => 211, b => 215, p => False), (a => 219, b => 223, p => False), (a => 227, b => 231, p => False), (a => 235, b => 239, p => False), (a => 243, b => 247, p => False), (a => 251, b => 255, p => False), (a => 259, b => 263, p => False), (a => 267, b => 271, p => False), (a => 275, b => 279, p => False), (a => 283, b => 287, p => False), (a => 291, b => 295, p => False), (a => 299, b => 303, p => False), (a => 307, b => 311, p => False), (a => 315, b => 319, p => False), (a => 323, b => 327, p => False), (a => 331, b => 335, p => False), (a => 339, b => 343, p => False), (a => 347, b => 351, p => False), (a => 66 , b => 70 , p => False), (a => 74 , b => 78 , p => False), (a => 82 , b => 86 , p => False), (a => 90 , b => 94 , p => False), (a => 98 , b => 102, p => False), (a => 106, b => 110, p => False), (a => 114, b => 118, p => False), (a => 122, b => 126, p => False), (a => 130, b => 134, p => False), (a => 138, b => 142, p => False), (a => 146, b => 150, p => False), (a => 154, b => 158, p => False), (a => 162, b => 166, p => False), (a => 170, b => 174, p => False), (a => 178, b => 182, p => False), (a => 186, b => 190, p => False), (a => 194, b => 198, p => False), (a => 202, b => 206, p => False), (a => 210, b => 214, p => False), (a => 218, b => 222, p => False), (a => 226, b => 230, p => False), (a => 234, b => 238, p => False), (a => 242, b => 246, p => False), (a => 250, b => 254, p => False), (a => 258, b => 262, p => False), (a => 266, b => 270, p => False), (a => 274, b => 278, p => False), (a => 282, b => 286, p => False), (a => 290, b => 294, p => False), (a => 298, b => 302, p => False), (a => 306, b => 310, p => False), (a => 314, b => 318, p => False), (a => 322, b => 326, p => False), (a => 330, b => 334, p => False), (a => 338, b => 342, p => False), (a => 346, b => 350, p => False), (a => 65 , b => 69 , p => False), (a => 73 , b => 77 , p => False), (a => 81 , b => 85 , p => False), (a => 89 , b => 93 , p => False), (a => 97 , b => 101, p => False), (a => 105, b => 109, p => False), (a => 113, b => 117, p => False), (a => 121, b => 125, p => False), (a => 129, b => 133, p => False), (a => 137, b => 141, p => False), (a => 145, b => 149, p => False), (a => 153, b => 157, p => False), (a => 161, b => 165, p => False), (a => 169, b => 173, p => False), (a => 177, b => 181, p => False), (a => 185, b => 189, p => False), (a => 193, b => 197, p => False), (a => 201, b => 205, p => False), (a => 209, b => 213, p => False), (a => 217, b => 221, p => False), (a => 225, b => 229, p => False), (a => 233, b => 237, p => False), (a => 241, b => 245, p => False), (a => 249, b => 253, p => False), (a => 257, b => 261, p => False), (a => 265, b => 269, p => False), (a => 273, b => 277, p => False), (a => 281, b => 285, p => False), (a => 289, b => 293, p => False), (a => 297, b => 301, p => False), (a => 305, b => 309, p => False), (a => 313, b => 317, p => False), (a => 321, b => 325, p => False), (a => 329, b => 333, p => False), (a => 337, b => 341, p => False), (a => 345, b => 349, p => False)),
                    ((a => 1  , b => 2  , p => False), (a => 5  , b => 6  , p => False), (a => 9  , b => 10 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 21 , b => 22 , p => False), (a => 25 , b => 26 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 37 , b => 38 , p => False), (a => 41 , b => 42 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 53 , b => 54 , p => False), (a => 57 , b => 58 , p => False), (a => 61 , b => 62 , p => False), (a => 0  , b => 4  , p => False), (a => 8  , b => 12 , p => False), (a => 16 , b => 20 , p => False), (a => 24 , b => 28 , p => False), (a => 32 , b => 36 , p => False), (a => 40 , b => 44 , p => False), (a => 48 , b => 52 , p => False), (a => 56 , b => 60 , p => False), (a => 3  , b => 7  , p => False), (a => 11 , b => 15 , p => False), (a => 19 , b => 23 , p => False), (a => 27 , b => 31 , p => False), (a => 35 , b => 39 , p => False), (a => 43 , b => 47 , p => False), (a => 51 , b => 55 , p => False), (a => 59 , b => 63 , p => False), (a => 64 , b => 72 , p => False), (a => 80 , b => 88 , p => False), (a => 96 , b => 104, p => False), (a => 112, b => 120, p => False), (a => 128, b => 136, p => False), (a => 144, b => 152, p => False), (a => 160, b => 168, p => False), (a => 176, b => 184, p => False), (a => 192, b => 200, p => False), (a => 208, b => 216, p => False), (a => 224, b => 232, p => False), (a => 240, b => 248, p => False), (a => 256, b => 264, p => False), (a => 272, b => 280, p => False), (a => 288, b => 296, p => False), (a => 304, b => 312, p => False), (a => 320, b => 328, p => False), (a => 336, b => 344, p => False), (a => 71 , b => 79 , p => False), (a => 87 , b => 95 , p => False), (a => 103, b => 111, p => False), (a => 119, b => 127, p => False), (a => 135, b => 143, p => False), (a => 151, b => 159, p => False), (a => 167, b => 175, p => False), (a => 183, b => 191, p => False), (a => 199, b => 207, p => False), (a => 215, b => 223, p => False), (a => 231, b => 239, p => False), (a => 247, b => 255, p => False), (a => 263, b => 271, p => False), (a => 279, b => 287, p => False), (a => 295, b => 303, p => False), (a => 311, b => 319, p => False), (a => 327, b => 335, p => False), (a => 343, b => 351, p => False), (a => 66 , b => 68 , p => False), (a => 74 , b => 76 , p => False), (a => 82 , b => 84 , p => False), (a => 90 , b => 92 , p => False), (a => 98 , b => 100, p => False), (a => 106, b => 108, p => False), (a => 114, b => 116, p => False), (a => 122, b => 124, p => False), (a => 130, b => 132, p => False), (a => 138, b => 140, p => False), (a => 146, b => 148, p => False), (a => 154, b => 156, p => False), (a => 162, b => 164, p => False), (a => 170, b => 172, p => False), (a => 178, b => 180, p => False), (a => 186, b => 188, p => False), (a => 194, b => 196, p => False), (a => 202, b => 204, p => False), (a => 210, b => 212, p => False), (a => 218, b => 220, p => False), (a => 226, b => 228, p => False), (a => 234, b => 236, p => False), (a => 242, b => 244, p => False), (a => 250, b => 252, p => False), (a => 258, b => 260, p => False), (a => 266, b => 268, p => False), (a => 274, b => 276, p => False), (a => 282, b => 284, p => False), (a => 290, b => 292, p => False), (a => 298, b => 300, p => False), (a => 306, b => 308, p => False), (a => 314, b => 316, p => False), (a => 322, b => 324, p => False), (a => 330, b => 332, p => False), (a => 338, b => 340, p => False), (a => 346, b => 348, p => False), (a => 67 , b => 69 , p => False), (a => 75 , b => 77 , p => False), (a => 83 , b => 85 , p => False), (a => 91 , b => 93 , p => False), (a => 99 , b => 101, p => False), (a => 107, b => 109, p => False), (a => 115, b => 117, p => False), (a => 123, b => 125, p => False), (a => 131, b => 133, p => False), (a => 139, b => 141, p => False), (a => 147, b => 149, p => False), (a => 155, b => 157, p => False), (a => 163, b => 165, p => False), (a => 171, b => 173, p => False), (a => 179, b => 181, p => False), (a => 187, b => 189, p => False), (a => 195, b => 197, p => False), (a => 203, b => 205, p => False), (a => 211, b => 213, p => False), (a => 219, b => 221, p => False), (a => 227, b => 229, p => False), (a => 235, b => 237, p => False), (a => 243, b => 245, p => False), (a => 251, b => 253, p => False), (a => 259, b => 261, p => False), (a => 267, b => 269, p => False), (a => 275, b => 277, p => False), (a => 283, b => 285, p => False), (a => 291, b => 293, p => False), (a => 299, b => 301, p => False), (a => 307, b => 309, p => False), (a => 315, b => 317, p => False), (a => 323, b => 325, p => False), (a => 331, b => 333, p => False), (a => 339, b => 341, p => False), (a => 347, b => 349, p => False), (a => 65 , b => 350, p => True ), (a => 70 , b => 345, p => True ), (a => 73 , b => 342, p => True ), (a => 78 , b => 337, p => True ), (a => 81 , b => 334, p => True ), (a => 86 , b => 329, p => True ), (a => 89 , b => 326, p => True ), (a => 94 , b => 321, p => True ), (a => 97 , b => 318, p => True ), (a => 102, b => 313, p => True ), (a => 105, b => 310, p => True ), (a => 110, b => 305, p => True ), (a => 113, b => 302, p => True ), (a => 118, b => 297, p => True ), (a => 121, b => 294, p => True ), (a => 126, b => 289, p => True ), (a => 129, b => 286, p => True ), (a => 134, b => 281, p => True ), (a => 137, b => 278, p => True ), (a => 142, b => 273, p => True ), (a => 145, b => 270, p => True ), (a => 150, b => 265, p => True ), (a => 153, b => 262, p => True ), (a => 158, b => 257, p => True ), (a => 161, b => 254, p => True ), (a => 166, b => 249, p => True ), (a => 169, b => 246, p => True ), (a => 174, b => 241, p => True ), (a => 177, b => 238, p => True ), (a => 182, b => 233, p => True ), (a => 185, b => 230, p => True ), (a => 190, b => 225, p => True ), (a => 193, b => 222, p => True ), (a => 198, b => 217, p => True ), (a => 201, b => 214, p => True ), (a => 206, b => 209, p => True )),
                    ((a => 2  , b => 6  , p => False), (a => 10 , b => 14 , p => False), (a => 18 , b => 22 , p => False), (a => 26 , b => 30 , p => False), (a => 34 , b => 38 , p => False), (a => 42 , b => 46 , p => False), (a => 50 , b => 54 , p => False), (a => 58 , b => 62 , p => False), (a => 1  , b => 5  , p => False), (a => 9  , b => 13 , p => False), (a => 17 , b => 21 , p => False), (a => 25 , b => 29 , p => False), (a => 33 , b => 37 , p => False), (a => 41 , b => 45 , p => False), (a => 49 , b => 53 , p => False), (a => 57 , b => 61 , p => False), (a => 0  , b => 8  , p => False), (a => 16 , b => 24 , p => False), (a => 32 , b => 40 , p => False), (a => 48 , b => 56 , p => False), (a => 7  , b => 15 , p => False), (a => 23 , b => 31 , p => False), (a => 39 , b => 47 , p => False), (a => 55 , b => 63 , p => False), (a => 64 , b => 80 , p => False), (a => 96 , b => 112, p => False), (a => 128, b => 144, p => False), (a => 160, b => 176, p => False), (a => 192, b => 208, p => False), (a => 224, b => 240, p => False), (a => 256, b => 272, p => False), (a => 288, b => 304, p => False), (a => 320, b => 336, p => False), (a => 79 , b => 95 , p => False), (a => 111, b => 127, p => False), (a => 143, b => 159, p => False), (a => 175, b => 191, p => False), (a => 207, b => 223, p => False), (a => 239, b => 255, p => False), (a => 271, b => 287, p => False), (a => 303, b => 319, p => False), (a => 335, b => 351, p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 89 , b => 90 , p => False), (a => 91 , b => 92 , p => False), (a => 93 , b => 94 , p => False), (a => 97 , b => 98 , p => False), (a => 99 , b => 100, p => False), (a => 101, b => 102, p => False), (a => 105, b => 106, p => False), (a => 107, b => 108, p => False), (a => 109, b => 110, p => False), (a => 113, b => 114, p => False), (a => 115, b => 116, p => False), (a => 117, b => 118, p => False), (a => 121, b => 122, p => False), (a => 123, b => 124, p => False), (a => 125, b => 126, p => False), (a => 129, b => 130, p => False), (a => 131, b => 132, p => False), (a => 133, b => 134, p => False), (a => 137, b => 138, p => False), (a => 139, b => 140, p => False), (a => 141, b => 142, p => False), (a => 145, b => 146, p => False), (a => 147, b => 148, p => False), (a => 149, b => 150, p => False), (a => 153, b => 154, p => False), (a => 155, b => 156, p => False), (a => 157, b => 158, p => False), (a => 161, b => 162, p => False), (a => 163, b => 164, p => False), (a => 165, b => 166, p => False), (a => 169, b => 170, p => False), (a => 171, b => 172, p => False), (a => 173, b => 174, p => False), (a => 177, b => 178, p => False), (a => 179, b => 180, p => False), (a => 181, b => 182, p => False), (a => 185, b => 186, p => False), (a => 187, b => 188, p => False), (a => 189, b => 190, p => False), (a => 193, b => 194, p => False), (a => 195, b => 196, p => False), (a => 197, b => 198, p => False), (a => 201, b => 202, p => False), (a => 203, b => 204, p => False), (a => 205, b => 206, p => False), (a => 209, b => 210, p => False), (a => 211, b => 212, p => False), (a => 213, b => 214, p => False), (a => 217, b => 218, p => False), (a => 219, b => 220, p => False), (a => 221, b => 222, p => False), (a => 225, b => 226, p => False), (a => 227, b => 228, p => False), (a => 229, b => 230, p => False), (a => 233, b => 234, p => False), (a => 235, b => 236, p => False), (a => 237, b => 238, p => False), (a => 241, b => 242, p => False), (a => 243, b => 244, p => False), (a => 245, b => 246, p => False), (a => 249, b => 250, p => False), (a => 251, b => 252, p => False), (a => 253, b => 254, p => False), (a => 257, b => 258, p => False), (a => 259, b => 260, p => False), (a => 261, b => 262, p => False), (a => 265, b => 266, p => False), (a => 267, b => 268, p => False), (a => 269, b => 270, p => False), (a => 273, b => 274, p => False), (a => 275, b => 276, p => False), (a => 277, b => 278, p => False), (a => 281, b => 282, p => False), (a => 283, b => 284, p => False), (a => 285, b => 286, p => False), (a => 289, b => 290, p => False), (a => 291, b => 292, p => False), (a => 293, b => 294, p => False), (a => 297, b => 298, p => False), (a => 299, b => 300, p => False), (a => 301, b => 302, p => False), (a => 305, b => 306, p => False), (a => 307, b => 308, p => False), (a => 309, b => 310, p => False), (a => 313, b => 314, p => False), (a => 315, b => 316, p => False), (a => 317, b => 318, p => False), (a => 321, b => 322, p => False), (a => 323, b => 324, p => False), (a => 325, b => 326, p => False), (a => 329, b => 330, p => False), (a => 331, b => 332, p => False), (a => 333, b => 334, p => False), (a => 337, b => 338, p => False), (a => 339, b => 340, p => False), (a => 341, b => 342, p => False), (a => 345, b => 346, p => False), (a => 347, b => 348, p => False), (a => 349, b => 350, p => False), (a => 3  , b => 344, p => True ), (a => 4  , b => 343, p => True ), (a => 11 , b => 328, p => True ), (a => 12 , b => 327, p => True ), (a => 19 , b => 312, p => True ), (a => 20 , b => 311, p => True ), (a => 27 , b => 296, p => True ), (a => 28 , b => 295, p => True ), (a => 35 , b => 280, p => True ), (a => 36 , b => 279, p => True ), (a => 43 , b => 264, p => True ), (a => 44 , b => 263, p => True ), (a => 51 , b => 248, p => True ), (a => 52 , b => 247, p => True ), (a => 59 , b => 232, p => True ), (a => 60 , b => 231, p => True ), (a => 71 , b => 216, p => True ), (a => 72 , b => 215, p => True ), (a => 87 , b => 200, p => True ), (a => 88 , b => 199, p => True ), (a => 103, b => 184, p => True ), (a => 104, b => 183, p => True ), (a => 119, b => 168, p => True ), (a => 120, b => 167, p => True ), (a => 135, b => 152, p => True ), (a => 136, b => 151, p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 10 , b => 12 , p => False), (a => 18 , b => 20 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 42 , b => 44 , p => False), (a => 50 , b => 52 , p => False), (a => 58 , b => 60 , p => False), (a => 3  , b => 5  , p => False), (a => 11 , b => 13 , p => False), (a => 19 , b => 21 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 43 , b => 45 , p => False), (a => 51 , b => 53 , p => False), (a => 59 , b => 61 , p => False), (a => 0  , b => 16 , p => False), (a => 32 , b => 48 , p => False), (a => 15 , b => 31 , p => False), (a => 47 , b => 63 , p => False), (a => 64 , b => 96 , p => False), (a => 128, b => 160, p => False), (a => 192, b => 224, p => False), (a => 256, b => 288, p => False), (a => 95 , b => 127, p => False), (a => 159, b => 191, p => False), (a => 223, b => 255, p => False), (a => 287, b => 319, p => False), (a => 68 , b => 76 , p => False), (a => 84 , b => 92 , p => False), (a => 100, b => 108, p => False), (a => 116, b => 124, p => False), (a => 132, b => 140, p => False), (a => 148, b => 156, p => False), (a => 164, b => 172, p => False), (a => 180, b => 188, p => False), (a => 196, b => 204, p => False), (a => 212, b => 220, p => False), (a => 228, b => 236, p => False), (a => 244, b => 252, p => False), (a => 260, b => 268, p => False), (a => 276, b => 284, p => False), (a => 292, b => 300, p => False), (a => 308, b => 316, p => False), (a => 324, b => 332, p => False), (a => 340, b => 348, p => False), (a => 66 , b => 74 , p => False), (a => 82 , b => 90 , p => False), (a => 98 , b => 106, p => False), (a => 114, b => 122, p => False), (a => 130, b => 138, p => False), (a => 146, b => 154, p => False), (a => 162, b => 170, p => False), (a => 178, b => 186, p => False), (a => 194, b => 202, p => False), (a => 210, b => 218, p => False), (a => 226, b => 234, p => False), (a => 242, b => 250, p => False), (a => 258, b => 266, p => False), (a => 274, b => 282, p => False), (a => 290, b => 298, p => False), (a => 306, b => 314, p => False), (a => 322, b => 330, p => False), (a => 338, b => 346, p => False), (a => 70 , b => 78 , p => False), (a => 86 , b => 94 , p => False), (a => 102, b => 110, p => False), (a => 118, b => 126, p => False), (a => 134, b => 142, p => False), (a => 150, b => 158, p => False), (a => 166, b => 174, p => False), (a => 182, b => 190, p => False), (a => 198, b => 206, p => False), (a => 214, b => 222, p => False), (a => 230, b => 238, p => False), (a => 246, b => 254, p => False), (a => 262, b => 270, p => False), (a => 278, b => 286, p => False), (a => 294, b => 302, p => False), (a => 310, b => 318, p => False), (a => 326, b => 334, p => False), (a => 342, b => 350, p => False), (a => 65 , b => 73 , p => False), (a => 81 , b => 89 , p => False), (a => 97 , b => 105, p => False), (a => 113, b => 121, p => False), (a => 129, b => 137, p => False), (a => 145, b => 153, p => False), (a => 161, b => 169, p => False), (a => 177, b => 185, p => False), (a => 193, b => 201, p => False), (a => 209, b => 217, p => False), (a => 225, b => 233, p => False), (a => 241, b => 249, p => False), (a => 257, b => 265, p => False), (a => 273, b => 281, p => False), (a => 289, b => 297, p => False), (a => 305, b => 313, p => False), (a => 321, b => 329, p => False), (a => 337, b => 345, p => False), (a => 69 , b => 77 , p => False), (a => 85 , b => 93 , p => False), (a => 101, b => 109, p => False), (a => 117, b => 125, p => False), (a => 133, b => 141, p => False), (a => 149, b => 157, p => False), (a => 165, b => 173, p => False), (a => 181, b => 189, p => False), (a => 197, b => 205, p => False), (a => 213, b => 221, p => False), (a => 229, b => 237, p => False), (a => 245, b => 253, p => False), (a => 261, b => 269, p => False), (a => 277, b => 285, p => False), (a => 293, b => 301, p => False), (a => 309, b => 317, p => False), (a => 325, b => 333, p => False), (a => 341, b => 349, p => False), (a => 67 , b => 75 , p => False), (a => 83 , b => 91 , p => False), (a => 99 , b => 107, p => False), (a => 115, b => 123, p => False), (a => 131, b => 139, p => False), (a => 147, b => 155, p => False), (a => 163, b => 171, p => False), (a => 179, b => 187, p => False), (a => 195, b => 203, p => False), (a => 211, b => 219, p => False), (a => 227, b => 235, p => False), (a => 243, b => 251, p => False), (a => 259, b => 267, p => False), (a => 275, b => 283, p => False), (a => 291, b => 299, p => False), (a => 307, b => 315, p => False), (a => 323, b => 331, p => False), (a => 339, b => 347, p => False), (a => 1  , b => 351, p => True ), (a => 6  , b => 344, p => True ), (a => 7  , b => 343, p => True ), (a => 8  , b => 336, p => True ), (a => 9  , b => 335, p => True ), (a => 14 , b => 328, p => True ), (a => 17 , b => 327, p => True ), (a => 22 , b => 320, p => True ), (a => 23 , b => 312, p => True ), (a => 24 , b => 311, p => True ), (a => 25 , b => 304, p => True ), (a => 30 , b => 303, p => True ), (a => 33 , b => 296, p => True ), (a => 38 , b => 295, p => True ), (a => 39 , b => 280, p => True ), (a => 40 , b => 279, p => True ), (a => 41 , b => 272, p => True ), (a => 46 , b => 271, p => True ), (a => 49 , b => 264, p => True ), (a => 54 , b => 263, p => True ), (a => 55 , b => 248, p => True ), (a => 56 , b => 247, p => True ), (a => 57 , b => 240, p => True ), (a => 62 , b => 239, p => True ), (a => 71 , b => 232, p => True ), (a => 72 , b => 231, p => True ), (a => 79 , b => 216, p => True ), (a => 80 , b => 215, p => True ), (a => 87 , b => 208, p => True ), (a => 88 , b => 207, p => True ), (a => 103, b => 200, p => True ), (a => 104, b => 199, p => True ), (a => 111, b => 184, p => True ), (a => 112, b => 183, p => True ), (a => 119, b => 176, p => True ), (a => 120, b => 175, p => True ), (a => 135, b => 168, p => True ), (a => 136, b => 167, p => True ), (a => 143, b => 152, p => True ), (a => 144, b => 151, p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 0  , b => 32 , p => False), (a => 31 , b => 63 , p => False), (a => 128, b => 192, p => False), (a => 256, b => 320, p => False), (a => 191, b => 255, p => False), (a => 68 , b => 72 , p => False), (a => 84 , b => 88 , p => False), (a => 100, b => 104, p => False), (a => 116, b => 120, p => False), (a => 132, b => 136, p => False), (a => 148, b => 152, p => False), (a => 164, b => 168, p => False), (a => 180, b => 184, p => False), (a => 196, b => 200, p => False), (a => 212, b => 216, p => False), (a => 228, b => 232, p => False), (a => 244, b => 248, p => False), (a => 260, b => 264, p => False), (a => 276, b => 280, p => False), (a => 292, b => 296, p => False), (a => 308, b => 312, p => False), (a => 324, b => 328, p => False), (a => 340, b => 344, p => False), (a => 70 , b => 74 , p => False), (a => 86 , b => 90 , p => False), (a => 102, b => 106, p => False), (a => 118, b => 122, p => False), (a => 134, b => 138, p => False), (a => 150, b => 154, p => False), (a => 166, b => 170, p => False), (a => 182, b => 186, p => False), (a => 198, b => 202, p => False), (a => 214, b => 218, p => False), (a => 230, b => 234, p => False), (a => 246, b => 250, p => False), (a => 262, b => 266, p => False), (a => 278, b => 282, p => False), (a => 294, b => 298, p => False), (a => 310, b => 314, p => False), (a => 326, b => 330, p => False), (a => 342, b => 346, p => False), (a => 69 , b => 73 , p => False), (a => 85 , b => 89 , p => False), (a => 101, b => 105, p => False), (a => 117, b => 121, p => False), (a => 133, b => 137, p => False), (a => 149, b => 153, p => False), (a => 165, b => 169, p => False), (a => 181, b => 185, p => False), (a => 197, b => 201, p => False), (a => 213, b => 217, p => False), (a => 229, b => 233, p => False), (a => 245, b => 249, p => False), (a => 261, b => 265, p => False), (a => 277, b => 281, p => False), (a => 293, b => 297, p => False), (a => 309, b => 313, p => False), (a => 325, b => 329, p => False), (a => 341, b => 345, p => False), (a => 71 , b => 75 , p => False), (a => 87 , b => 91 , p => False), (a => 103, b => 107, p => False), (a => 119, b => 123, p => False), (a => 135, b => 139, p => False), (a => 151, b => 155, p => False), (a => 167, b => 171, p => False), (a => 183, b => 187, p => False), (a => 199, b => 203, p => False), (a => 215, b => 219, p => False), (a => 231, b => 235, p => False), (a => 247, b => 251, p => False), (a => 263, b => 267, p => False), (a => 279, b => 283, p => False), (a => 295, b => 299, p => False), (a => 311, b => 315, p => False), (a => 327, b => 331, p => False), (a => 343, b => 347, p => False), (a => 7  , b => 351, p => True ), (a => 8  , b => 350, p => True ), (a => 15 , b => 349, p => True ), (a => 16 , b => 348, p => True ), (a => 23 , b => 339, p => True ), (a => 24 , b => 338, p => True ), (a => 39 , b => 337, p => True ), (a => 40 , b => 336, p => True ), (a => 47 , b => 335, p => True ), (a => 48 , b => 334, p => True ), (a => 55 , b => 333, p => True ), (a => 56 , b => 332, p => True ), (a => 64 , b => 323, p => True ), (a => 65 , b => 322, p => True ), (a => 66 , b => 321, p => True ), (a => 67 , b => 319, p => True ), (a => 76 , b => 318, p => True ), (a => 77 , b => 317, p => True ), (a => 78 , b => 316, p => True ), (a => 79 , b => 307, p => True ), (a => 80 , b => 306, p => True ), (a => 81 , b => 305, p => True ), (a => 82 , b => 304, p => True ), (a => 83 , b => 303, p => True ), (a => 92 , b => 302, p => True ), (a => 93 , b => 301, p => True ), (a => 94 , b => 300, p => True ), (a => 95 , b => 291, p => True ), (a => 96 , b => 290, p => True ), (a => 97 , b => 289, p => True ), (a => 98 , b => 288, p => True ), (a => 99 , b => 287, p => True ), (a => 108, b => 286, p => True ), (a => 109, b => 285, p => True ), (a => 110, b => 284, p => True ), (a => 111, b => 275, p => True ), (a => 112, b => 274, p => True ), (a => 113, b => 273, p => True ), (a => 114, b => 272, p => True ), (a => 115, b => 271, p => True ), (a => 124, b => 270, p => True ), (a => 125, b => 269, p => True ), (a => 126, b => 268, p => True ), (a => 127, b => 259, p => True ), (a => 129, b => 258, p => True ), (a => 130, b => 257, p => True ), (a => 131, b => 254, p => True ), (a => 140, b => 253, p => True ), (a => 141, b => 252, p => True ), (a => 142, b => 243, p => True ), (a => 143, b => 242, p => True ), (a => 144, b => 241, p => True ), (a => 145, b => 240, p => True ), (a => 146, b => 239, p => True ), (a => 147, b => 238, p => True ), (a => 156, b => 237, p => True ), (a => 157, b => 236, p => True ), (a => 158, b => 227, p => True ), (a => 159, b => 226, p => True ), (a => 160, b => 225, p => True ), (a => 161, b => 224, p => True ), (a => 162, b => 223, p => True ), (a => 163, b => 222, p => True ), (a => 172, b => 221, p => True ), (a => 173, b => 220, p => True ), (a => 174, b => 211, p => True ), (a => 175, b => 210, p => True ), (a => 176, b => 209, p => True ), (a => 177, b => 208, p => True ), (a => 178, b => 207, p => True ), (a => 179, b => 206, p => True ), (a => 188, b => 205, p => True ), (a => 189, b => 204, p => True ), (a => 190, b => 195, p => True ), (a => 193, b => 194, p => True )),
                    ((a => 4  , b => 12 , p => False), (a => 20 , b => 28 , p => False), (a => 36 , b => 44 , p => False), (a => 52 , b => 60 , p => False), (a => 2  , b => 10 , p => False), (a => 18 , b => 26 , p => False), (a => 34 , b => 42 , p => False), (a => 50 , b => 58 , p => False), (a => 6  , b => 14 , p => False), (a => 22 , b => 30 , p => False), (a => 38 , b => 46 , p => False), (a => 54 , b => 62 , p => False), (a => 1  , b => 9  , p => False), (a => 17 , b => 25 , p => False), (a => 33 , b => 41 , p => False), (a => 49 , b => 57 , p => False), (a => 5  , b => 13 , p => False), (a => 21 , b => 29 , p => False), (a => 37 , b => 45 , p => False), (a => 53 , b => 61 , p => False), (a => 3  , b => 11 , p => False), (a => 19 , b => 27 , p => False), (a => 35 , b => 43 , p => False), (a => 51 , b => 59 , p => False), (a => 0  , b => 64 , p => False), (a => 63 , b => 127, p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 82 , b => 84 , p => False), (a => 86 , b => 88 , p => False), (a => 90 , b => 92 , p => False), (a => 98 , b => 100, p => False), (a => 102, b => 104, p => False), (a => 106, b => 108, p => False), (a => 114, b => 116, p => False), (a => 118, b => 120, p => False), (a => 122, b => 124, p => False), (a => 130, b => 132, p => False), (a => 134, b => 136, p => False), (a => 138, b => 140, p => False), (a => 146, b => 148, p => False), (a => 150, b => 152, p => False), (a => 154, b => 156, p => False), (a => 162, b => 164, p => False), (a => 166, b => 168, p => False), (a => 170, b => 172, p => False), (a => 178, b => 180, p => False), (a => 182, b => 184, p => False), (a => 186, b => 188, p => False), (a => 194, b => 196, p => False), (a => 198, b => 200, p => False), (a => 202, b => 204, p => False), (a => 210, b => 212, p => False), (a => 214, b => 216, p => False), (a => 218, b => 220, p => False), (a => 226, b => 228, p => False), (a => 230, b => 232, p => False), (a => 234, b => 236, p => False), (a => 242, b => 244, p => False), (a => 246, b => 248, p => False), (a => 250, b => 252, p => False), (a => 258, b => 260, p => False), (a => 262, b => 264, p => False), (a => 266, b => 268, p => False), (a => 274, b => 276, p => False), (a => 278, b => 280, p => False), (a => 282, b => 284, p => False), (a => 290, b => 292, p => False), (a => 294, b => 296, p => False), (a => 298, b => 300, p => False), (a => 306, b => 308, p => False), (a => 310, b => 312, p => False), (a => 314, b => 316, p => False), (a => 322, b => 324, p => False), (a => 326, b => 328, p => False), (a => 330, b => 332, p => False), (a => 338, b => 340, p => False), (a => 342, b => 344, p => False), (a => 346, b => 348, p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 83 , b => 85 , p => False), (a => 87 , b => 89 , p => False), (a => 91 , b => 93 , p => False), (a => 99 , b => 101, p => False), (a => 103, b => 105, p => False), (a => 107, b => 109, p => False), (a => 115, b => 117, p => False), (a => 119, b => 121, p => False), (a => 123, b => 125, p => False), (a => 131, b => 133, p => False), (a => 135, b => 137, p => False), (a => 139, b => 141, p => False), (a => 147, b => 149, p => False), (a => 151, b => 153, p => False), (a => 155, b => 157, p => False), (a => 163, b => 165, p => False), (a => 167, b => 169, p => False), (a => 171, b => 173, p => False), (a => 179, b => 181, p => False), (a => 183, b => 185, p => False), (a => 187, b => 189, p => False), (a => 195, b => 197, p => False), (a => 199, b => 201, p => False), (a => 203, b => 205, p => False), (a => 211, b => 213, p => False), (a => 215, b => 217, p => False), (a => 219, b => 221, p => False), (a => 227, b => 229, p => False), (a => 231, b => 233, p => False), (a => 235, b => 237, p => False), (a => 243, b => 245, p => False), (a => 247, b => 249, p => False), (a => 251, b => 253, p => False), (a => 259, b => 261, p => False), (a => 263, b => 265, p => False), (a => 267, b => 269, p => False), (a => 275, b => 277, p => False), (a => 279, b => 281, p => False), (a => 283, b => 285, p => False), (a => 291, b => 293, p => False), (a => 295, b => 297, p => False), (a => 299, b => 301, p => False), (a => 307, b => 309, p => False), (a => 311, b => 313, p => False), (a => 315, b => 317, p => False), (a => 323, b => 325, p => False), (a => 327, b => 329, p => False), (a => 331, b => 333, p => False), (a => 339, b => 341, p => False), (a => 343, b => 345, p => False), (a => 347, b => 349, p => False), (a => 7  , b => 351, p => True ), (a => 8  , b => 350, p => True ), (a => 15 , b => 337, p => True ), (a => 16 , b => 336, p => True ), (a => 23 , b => 335, p => True ), (a => 24 , b => 334, p => True ), (a => 31 , b => 321, p => True ), (a => 32 , b => 320, p => True ), (a => 39 , b => 319, p => True ), (a => 40 , b => 318, p => True ), (a => 47 , b => 305, p => True ), (a => 48 , b => 304, p => True ), (a => 55 , b => 303, p => True ), (a => 56 , b => 302, p => True ), (a => 65 , b => 289, p => True ), (a => 78 , b => 288, p => True ), (a => 79 , b => 287, p => True ), (a => 80 , b => 286, p => True ), (a => 81 , b => 273, p => True ), (a => 94 , b => 272, p => True ), (a => 95 , b => 271, p => True ), (a => 96 , b => 270, p => True ), (a => 97 , b => 257, p => True ), (a => 110, b => 256, p => True ), (a => 111, b => 255, p => True ), (a => 112, b => 254, p => True ), (a => 113, b => 241, p => True ), (a => 126, b => 240, p => True ), (a => 128, b => 239, p => True ), (a => 129, b => 238, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 20 , b => 24 , p => False), (a => 36 , b => 40 , p => False), (a => 52 , b => 56 , p => False), (a => 6  , b => 10 , p => False), (a => 22 , b => 26 , p => False), (a => 38 , b => 42 , p => False), (a => 54 , b => 58 , p => False), (a => 5  , b => 9  , p => False), (a => 21 , b => 25 , p => False), (a => 37 , b => 41 , p => False), (a => 53 , b => 57 , p => False), (a => 7  , b => 11 , p => False), (a => 23 , b => 27 , p => False), (a => 39 , b => 43 , p => False), (a => 55 , b => 59 , p => False), (a => 0  , b => 128, p => False), (a => 127, b => 255, p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 87 , b => 88 , p => False), (a => 89 , b => 90 , p => False), (a => 91 , b => 92 , p => False), (a => 93 , b => 94 , p => False), (a => 97 , b => 98 , p => False), (a => 99 , b => 100, p => False), (a => 101, b => 102, p => False), (a => 103, b => 104, p => False), (a => 105, b => 106, p => False), (a => 107, b => 108, p => False), (a => 109, b => 110, p => False), (a => 113, b => 114, p => False), (a => 115, b => 116, p => False), (a => 117, b => 118, p => False), (a => 119, b => 120, p => False), (a => 121, b => 122, p => False), (a => 123, b => 124, p => False), (a => 125, b => 126, p => False), (a => 129, b => 130, p => False), (a => 131, b => 132, p => False), (a => 133, b => 134, p => False), (a => 135, b => 136, p => False), (a => 137, b => 138, p => False), (a => 139, b => 140, p => False), (a => 141, b => 142, p => False), (a => 145, b => 146, p => False), (a => 147, b => 148, p => False), (a => 149, b => 150, p => False), (a => 151, b => 152, p => False), (a => 153, b => 154, p => False), (a => 155, b => 156, p => False), (a => 157, b => 158, p => False), (a => 161, b => 162, p => False), (a => 163, b => 164, p => False), (a => 165, b => 166, p => False), (a => 167, b => 168, p => False), (a => 169, b => 170, p => False), (a => 171, b => 172, p => False), (a => 173, b => 174, p => False), (a => 177, b => 178, p => False), (a => 179, b => 180, p => False), (a => 181, b => 182, p => False), (a => 183, b => 184, p => False), (a => 185, b => 186, p => False), (a => 187, b => 188, p => False), (a => 189, b => 190, p => False), (a => 193, b => 194, p => False), (a => 195, b => 196, p => False), (a => 197, b => 198, p => False), (a => 199, b => 200, p => False), (a => 201, b => 202, p => False), (a => 203, b => 204, p => False), (a => 205, b => 206, p => False), (a => 209, b => 210, p => False), (a => 211, b => 212, p => False), (a => 213, b => 214, p => False), (a => 215, b => 216, p => False), (a => 217, b => 218, p => False), (a => 219, b => 220, p => False), (a => 221, b => 222, p => False), (a => 225, b => 226, p => False), (a => 227, b => 228, p => False), (a => 229, b => 230, p => False), (a => 231, b => 232, p => False), (a => 233, b => 234, p => False), (a => 235, b => 236, p => False), (a => 237, b => 238, p => False), (a => 241, b => 242, p => False), (a => 243, b => 244, p => False), (a => 245, b => 246, p => False), (a => 247, b => 248, p => False), (a => 249, b => 250, p => False), (a => 251, b => 252, p => False), (a => 253, b => 254, p => False), (a => 257, b => 258, p => False), (a => 259, b => 260, p => False), (a => 261, b => 262, p => False), (a => 263, b => 264, p => False), (a => 265, b => 266, p => False), (a => 267, b => 268, p => False), (a => 269, b => 270, p => False), (a => 273, b => 274, p => False), (a => 275, b => 276, p => False), (a => 277, b => 278, p => False), (a => 279, b => 280, p => False), (a => 281, b => 282, p => False), (a => 283, b => 284, p => False), (a => 285, b => 286, p => False), (a => 289, b => 290, p => False), (a => 291, b => 292, p => False), (a => 293, b => 294, p => False), (a => 295, b => 296, p => False), (a => 297, b => 298, p => False), (a => 299, b => 300, p => False), (a => 301, b => 302, p => False), (a => 305, b => 306, p => False), (a => 307, b => 308, p => False), (a => 309, b => 310, p => False), (a => 311, b => 312, p => False), (a => 313, b => 314, p => False), (a => 315, b => 316, p => False), (a => 317, b => 318, p => False), (a => 321, b => 322, p => False), (a => 323, b => 324, p => False), (a => 325, b => 326, p => False), (a => 327, b => 328, p => False), (a => 329, b => 330, p => False), (a => 331, b => 332, p => False), (a => 333, b => 334, p => False), (a => 337, b => 338, p => False), (a => 339, b => 340, p => False), (a => 341, b => 342, p => False), (a => 343, b => 344, p => False), (a => 345, b => 346, p => False), (a => 347, b => 348, p => False), (a => 349, b => 350, p => False), (a => 1  , b => 351, p => True ), (a => 2  , b => 336, p => True ), (a => 3  , b => 335, p => True ), (a => 12 , b => 320, p => True ), (a => 13 , b => 319, p => True ), (a => 14 , b => 304, p => True ), (a => 15 , b => 303, p => True ), (a => 16 , b => 288, p => True ), (a => 17 , b => 287, p => True ), (a => 18 , b => 272, p => True ), (a => 19 , b => 271, p => True ), (a => 28 , b => 256, p => True ), (a => 29 , b => 240, p => True ), (a => 30 , b => 239, p => True ), (a => 31 , b => 224, p => True ), (a => 32 , b => 223, p => True ), (a => 33 , b => 208, p => True ), (a => 34 , b => 207, p => True ), (a => 35 , b => 192, p => True ), (a => 44 , b => 191, p => True ), (a => 45 , b => 176, p => True ), (a => 46 , b => 175, p => True ), (a => 47 , b => 160, p => True ), (a => 48 , b => 159, p => True ), (a => 49 , b => 144, p => True ), (a => 50 , b => 143, p => True ), (a => 51 , b => 112, p => True ), (a => 60 , b => 111, p => True ), (a => 61 , b => 96 , p => True ), (a => 62 , b => 95 , p => True ), (a => 63 , b => 80 , p => True ), (a => 64 , b => 79 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 0  , b => 256, p => False), (a => 72 , b => 88 , p => False), (a => 104, b => 120, p => False), (a => 136, b => 152, p => False), (a => 168, b => 184, p => False), (a => 200, b => 216, p => False), (a => 232, b => 248, p => False), (a => 264, b => 280, p => False), (a => 296, b => 312, p => False), (a => 328, b => 344, p => False), (a => 68 , b => 84 , p => False), (a => 100, b => 116, p => False), (a => 132, b => 148, p => False), (a => 164, b => 180, p => False), (a => 196, b => 212, p => False), (a => 228, b => 244, p => False), (a => 260, b => 276, p => False), (a => 292, b => 308, p => False), (a => 324, b => 340, p => False), (a => 76 , b => 92 , p => False), (a => 108, b => 124, p => False), (a => 140, b => 156, p => False), (a => 172, b => 188, p => False), (a => 204, b => 220, p => False), (a => 236, b => 252, p => False), (a => 268, b => 284, p => False), (a => 300, b => 316, p => False), (a => 332, b => 348, p => False), (a => 66 , b => 82 , p => False), (a => 98 , b => 114, p => False), (a => 130, b => 146, p => False), (a => 162, b => 178, p => False), (a => 194, b => 210, p => False), (a => 226, b => 242, p => False), (a => 258, b => 274, p => False), (a => 290, b => 306, p => False), (a => 322, b => 338, p => False), (a => 74 , b => 90 , p => False), (a => 106, b => 122, p => False), (a => 138, b => 154, p => False), (a => 170, b => 186, p => False), (a => 202, b => 218, p => False), (a => 234, b => 250, p => False), (a => 266, b => 282, p => False), (a => 298, b => 314, p => False), (a => 330, b => 346, p => False), (a => 70 , b => 86 , p => False), (a => 102, b => 118, p => False), (a => 134, b => 150, p => False), (a => 166, b => 182, p => False), (a => 198, b => 214, p => False), (a => 230, b => 246, p => False), (a => 262, b => 278, p => False), (a => 294, b => 310, p => False), (a => 326, b => 342, p => False), (a => 78 , b => 94 , p => False), (a => 110, b => 126, p => False), (a => 142, b => 158, p => False), (a => 174, b => 190, p => False), (a => 206, b => 222, p => False), (a => 238, b => 254, p => False), (a => 270, b => 286, p => False), (a => 302, b => 318, p => False), (a => 334, b => 350, p => False), (a => 65 , b => 81 , p => False), (a => 97 , b => 113, p => False), (a => 129, b => 145, p => False), (a => 161, b => 177, p => False), (a => 193, b => 209, p => False), (a => 225, b => 241, p => False), (a => 257, b => 273, p => False), (a => 289, b => 305, p => False), (a => 321, b => 337, p => False), (a => 73 , b => 89 , p => False), (a => 105, b => 121, p => False), (a => 137, b => 153, p => False), (a => 169, b => 185, p => False), (a => 201, b => 217, p => False), (a => 233, b => 249, p => False), (a => 265, b => 281, p => False), (a => 297, b => 313, p => False), (a => 329, b => 345, p => False), (a => 69 , b => 85 , p => False), (a => 101, b => 117, p => False), (a => 133, b => 149, p => False), (a => 165, b => 181, p => False), (a => 197, b => 213, p => False), (a => 229, b => 245, p => False), (a => 261, b => 277, p => False), (a => 293, b => 309, p => False), (a => 325, b => 341, p => False), (a => 77 , b => 93 , p => False), (a => 109, b => 125, p => False), (a => 141, b => 157, p => False), (a => 173, b => 189, p => False), (a => 205, b => 221, p => False), (a => 237, b => 253, p => False), (a => 269, b => 285, p => False), (a => 301, b => 317, p => False), (a => 333, b => 349, p => False), (a => 67 , b => 83 , p => False), (a => 99 , b => 115, p => False), (a => 131, b => 147, p => False), (a => 163, b => 179, p => False), (a => 195, b => 211, p => False), (a => 227, b => 243, p => False), (a => 259, b => 275, p => False), (a => 291, b => 307, p => False), (a => 323, b => 339, p => False), (a => 75 , b => 91 , p => False), (a => 107, b => 123, p => False), (a => 139, b => 155, p => False), (a => 171, b => 187, p => False), (a => 203, b => 219, p => False), (a => 235, b => 251, p => False), (a => 267, b => 283, p => False), (a => 299, b => 315, p => False), (a => 331, b => 347, p => False), (a => 71 , b => 87 , p => False), (a => 103, b => 119, p => False), (a => 135, b => 151, p => False), (a => 167, b => 183, p => False), (a => 199, b => 215, p => False), (a => 231, b => 247, p => False), (a => 263, b => 279, p => False), (a => 295, b => 311, p => False), (a => 327, b => 343, p => False), (a => 1  , b => 351, p => True ), (a => 14 , b => 336, p => True ), (a => 15 , b => 335, p => True ), (a => 16 , b => 320, p => True ), (a => 17 , b => 319, p => True ), (a => 30 , b => 304, p => True ), (a => 31 , b => 303, p => True ), (a => 32 , b => 288, p => True ), (a => 33 , b => 287, p => True ), (a => 46 , b => 272, p => True ), (a => 47 , b => 271, p => True ), (a => 48 , b => 255, p => True ), (a => 49 , b => 240, p => True ), (a => 62 , b => 239, p => True ), (a => 63 , b => 224, p => True ), (a => 64 , b => 223, p => True ), (a => 79 , b => 208, p => True ), (a => 80 , b => 207, p => True ), (a => 95 , b => 192, p => True ), (a => 96 , b => 191, p => True ), (a => 111, b => 176, p => True ), (a => 112, b => 175, p => True ), (a => 127, b => 160, p => True ), (a => 128, b => 159, p => True ), (a => 143, b => 144, p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 72 , b => 80 , p => False), (a => 104, b => 112, p => False), (a => 136, b => 144, p => False), (a => 168, b => 176, p => False), (a => 200, b => 208, p => False), (a => 232, b => 240, p => False), (a => 264, b => 272, p => False), (a => 296, b => 304, p => False), (a => 328, b => 336, p => False), (a => 76 , b => 84 , p => False), (a => 108, b => 116, p => False), (a => 140, b => 148, p => False), (a => 172, b => 180, p => False), (a => 204, b => 212, p => False), (a => 236, b => 244, p => False), (a => 268, b => 276, p => False), (a => 300, b => 308, p => False), (a => 332, b => 340, p => False), (a => 74 , b => 82 , p => False), (a => 106, b => 114, p => False), (a => 138, b => 146, p => False), (a => 170, b => 178, p => False), (a => 202, b => 210, p => False), (a => 234, b => 242, p => False), (a => 266, b => 274, p => False), (a => 298, b => 306, p => False), (a => 330, b => 338, p => False), (a => 78 , b => 86 , p => False), (a => 110, b => 118, p => False), (a => 142, b => 150, p => False), (a => 174, b => 182, p => False), (a => 206, b => 214, p => False), (a => 238, b => 246, p => False), (a => 270, b => 278, p => False), (a => 302, b => 310, p => False), (a => 334, b => 342, p => False), (a => 73 , b => 81 , p => False), (a => 105, b => 113, p => False), (a => 137, b => 145, p => False), (a => 169, b => 177, p => False), (a => 201, b => 209, p => False), (a => 233, b => 241, p => False), (a => 265, b => 273, p => False), (a => 297, b => 305, p => False), (a => 329, b => 337, p => False), (a => 77 , b => 85 , p => False), (a => 109, b => 117, p => False), (a => 141, b => 149, p => False), (a => 173, b => 181, p => False), (a => 205, b => 213, p => False), (a => 237, b => 245, p => False), (a => 269, b => 277, p => False), (a => 301, b => 309, p => False), (a => 333, b => 341, p => False), (a => 75 , b => 83 , p => False), (a => 107, b => 115, p => False), (a => 139, b => 147, p => False), (a => 171, b => 179, p => False), (a => 203, b => 211, p => False), (a => 235, b => 243, p => False), (a => 267, b => 275, p => False), (a => 299, b => 307, p => False), (a => 331, b => 339, p => False), (a => 79 , b => 87 , p => False), (a => 111, b => 119, p => False), (a => 143, b => 151, p => False), (a => 175, b => 183, p => False), (a => 207, b => 215, p => False), (a => 239, b => 247, p => False), (a => 271, b => 279, p => False), (a => 303, b => 311, p => False), (a => 335, b => 343, p => False), (a => 0  , b => 351, p => True ), (a => 15 , b => 350, p => True ), (a => 16 , b => 349, p => True ), (a => 31 , b => 348, p => True ), (a => 32 , b => 347, p => True ), (a => 47 , b => 346, p => True ), (a => 48 , b => 345, p => True ), (a => 63 , b => 344, p => True ), (a => 64 , b => 327, p => True ), (a => 65 , b => 326, p => True ), (a => 66 , b => 325, p => True ), (a => 67 , b => 324, p => True ), (a => 68 , b => 323, p => True ), (a => 69 , b => 322, p => True ), (a => 70 , b => 321, p => True ), (a => 71 , b => 320, p => True ), (a => 88 , b => 319, p => True ), (a => 89 , b => 318, p => True ), (a => 90 , b => 317, p => True ), (a => 91 , b => 316, p => True ), (a => 92 , b => 315, p => True ), (a => 93 , b => 314, p => True ), (a => 94 , b => 313, p => True ), (a => 95 , b => 312, p => True ), (a => 96 , b => 295, p => True ), (a => 97 , b => 294, p => True ), (a => 98 , b => 293, p => True ), (a => 99 , b => 292, p => True ), (a => 100, b => 291, p => True ), (a => 101, b => 290, p => True ), (a => 102, b => 289, p => True ), (a => 103, b => 288, p => True ), (a => 120, b => 287, p => True ), (a => 121, b => 286, p => True ), (a => 122, b => 285, p => True ), (a => 123, b => 284, p => True ), (a => 124, b => 283, p => True ), (a => 125, b => 282, p => True ), (a => 126, b => 281, p => True ), (a => 127, b => 280, p => True ), (a => 128, b => 263, p => True ), (a => 129, b => 262, p => True ), (a => 130, b => 261, p => True ), (a => 131, b => 260, p => True ), (a => 132, b => 259, p => True ), (a => 133, b => 258, p => True ), (a => 134, b => 257, p => True ), (a => 135, b => 256, p => True ), (a => 152, b => 255, p => True ), (a => 153, b => 254, p => True ), (a => 154, b => 253, p => True ), (a => 155, b => 252, p => True ), (a => 156, b => 251, p => True ), (a => 157, b => 250, p => True ), (a => 158, b => 249, p => True ), (a => 159, b => 248, p => True ), (a => 160, b => 231, p => True ), (a => 161, b => 230, p => True ), (a => 162, b => 229, p => True ), (a => 163, b => 228, p => True ), (a => 164, b => 227, p => True ), (a => 165, b => 226, p => True ), (a => 166, b => 225, p => True ), (a => 167, b => 224, p => True ), (a => 184, b => 223, p => True ), (a => 185, b => 222, p => True ), (a => 186, b => 221, p => True ), (a => 187, b => 220, p => True ), (a => 188, b => 219, p => True ), (a => 189, b => 218, p => True ), (a => 190, b => 217, p => True ), (a => 191, b => 216, p => True ), (a => 192, b => 199, p => True ), (a => 193, b => 198, p => True ), (a => 194, b => 197, p => True ), (a => 195, b => 196, p => True )),
                    ((a => 8  , b => 24 , p => False), (a => 40 , b => 56 , p => False), (a => 4  , b => 20 , p => False), (a => 36 , b => 52 , p => False), (a => 12 , b => 28 , p => False), (a => 44 , b => 60 , p => False), (a => 2  , b => 18 , p => False), (a => 34 , b => 50 , p => False), (a => 10 , b => 26 , p => False), (a => 42 , b => 58 , p => False), (a => 6  , b => 22 , p => False), (a => 38 , b => 54 , p => False), (a => 14 , b => 30 , p => False), (a => 46 , b => 62 , p => False), (a => 1  , b => 17 , p => False), (a => 33 , b => 49 , p => False), (a => 9  , b => 25 , p => False), (a => 41 , b => 57 , p => False), (a => 5  , b => 21 , p => False), (a => 37 , b => 53 , p => False), (a => 13 , b => 29 , p => False), (a => 45 , b => 61 , p => False), (a => 3  , b => 19 , p => False), (a => 35 , b => 51 , p => False), (a => 11 , b => 27 , p => False), (a => 43 , b => 59 , p => False), (a => 7  , b => 23 , p => False), (a => 39 , b => 55 , p => False), (a => 68 , b => 72 , p => False), (a => 76 , b => 80 , p => False), (a => 84 , b => 88 , p => False), (a => 100, b => 104, p => False), (a => 108, b => 112, p => False), (a => 116, b => 120, p => False), (a => 132, b => 136, p => False), (a => 140, b => 144, p => False), (a => 148, b => 152, p => False), (a => 164, b => 168, p => False), (a => 172, b => 176, p => False), (a => 180, b => 184, p => False), (a => 196, b => 200, p => False), (a => 204, b => 208, p => False), (a => 212, b => 216, p => False), (a => 228, b => 232, p => False), (a => 236, b => 240, p => False), (a => 244, b => 248, p => False), (a => 260, b => 264, p => False), (a => 268, b => 272, p => False), (a => 276, b => 280, p => False), (a => 292, b => 296, p => False), (a => 300, b => 304, p => False), (a => 308, b => 312, p => False), (a => 324, b => 328, p => False), (a => 332, b => 336, p => False), (a => 340, b => 344, p => False), (a => 70 , b => 74 , p => False), (a => 78 , b => 82 , p => False), (a => 86 , b => 90 , p => False), (a => 102, b => 106, p => False), (a => 110, b => 114, p => False), (a => 118, b => 122, p => False), (a => 134, b => 138, p => False), (a => 142, b => 146, p => False), (a => 150, b => 154, p => False), (a => 166, b => 170, p => False), (a => 174, b => 178, p => False), (a => 182, b => 186, p => False), (a => 198, b => 202, p => False), (a => 206, b => 210, p => False), (a => 214, b => 218, p => False), (a => 230, b => 234, p => False), (a => 238, b => 242, p => False), (a => 246, b => 250, p => False), (a => 262, b => 266, p => False), (a => 270, b => 274, p => False), (a => 278, b => 282, p => False), (a => 294, b => 298, p => False), (a => 302, b => 306, p => False), (a => 310, b => 314, p => False), (a => 326, b => 330, p => False), (a => 334, b => 338, p => False), (a => 342, b => 346, p => False), (a => 69 , b => 73 , p => False), (a => 77 , b => 81 , p => False), (a => 85 , b => 89 , p => False), (a => 101, b => 105, p => False), (a => 109, b => 113, p => False), (a => 117, b => 121, p => False), (a => 133, b => 137, p => False), (a => 141, b => 145, p => False), (a => 149, b => 153, p => False), (a => 165, b => 169, p => False), (a => 173, b => 177, p => False), (a => 181, b => 185, p => False), (a => 197, b => 201, p => False), (a => 205, b => 209, p => False), (a => 213, b => 217, p => False), (a => 229, b => 233, p => False), (a => 237, b => 241, p => False), (a => 245, b => 249, p => False), (a => 261, b => 265, p => False), (a => 269, b => 273, p => False), (a => 277, b => 281, p => False), (a => 293, b => 297, p => False), (a => 301, b => 305, p => False), (a => 309, b => 313, p => False), (a => 325, b => 329, p => False), (a => 333, b => 337, p => False), (a => 341, b => 345, p => False), (a => 71 , b => 75 , p => False), (a => 79 , b => 83 , p => False), (a => 87 , b => 91 , p => False), (a => 103, b => 107, p => False), (a => 111, b => 115, p => False), (a => 119, b => 123, p => False), (a => 135, b => 139, p => False), (a => 143, b => 147, p => False), (a => 151, b => 155, p => False), (a => 167, b => 171, p => False), (a => 175, b => 179, p => False), (a => 183, b => 187, p => False), (a => 199, b => 203, p => False), (a => 207, b => 211, p => False), (a => 215, b => 219, p => False), (a => 231, b => 235, p => False), (a => 239, b => 243, p => False), (a => 247, b => 251, p => False), (a => 263, b => 267, p => False), (a => 271, b => 275, p => False), (a => 279, b => 283, p => False), (a => 295, b => 299, p => False), (a => 303, b => 307, p => False), (a => 311, b => 315, p => False), (a => 327, b => 331, p => False), (a => 335, b => 339, p => False), (a => 343, b => 347, p => False), (a => 0  , b => 351, p => True ), (a => 15 , b => 350, p => True ), (a => 16 , b => 349, p => True ), (a => 31 , b => 348, p => True ), (a => 32 , b => 323, p => True ), (a => 47 , b => 322, p => True ), (a => 48 , b => 321, p => True ), (a => 63 , b => 320, p => True ), (a => 64 , b => 319, p => True ), (a => 65 , b => 318, p => True ), (a => 66 , b => 317, p => True ), (a => 67 , b => 316, p => True ), (a => 92 , b => 291, p => True ), (a => 93 , b => 290, p => True ), (a => 94 , b => 289, p => True ), (a => 95 , b => 288, p => True ), (a => 96 , b => 287, p => True ), (a => 97 , b => 286, p => True ), (a => 98 , b => 285, p => True ), (a => 99 , b => 284, p => True ), (a => 124, b => 259, p => True ), (a => 125, b => 258, p => True ), (a => 126, b => 257, p => True ), (a => 127, b => 256, p => True ), (a => 128, b => 255, p => True ), (a => 129, b => 254, p => True ), (a => 130, b => 253, p => True ), (a => 131, b => 252, p => True ), (a => 156, b => 227, p => True ), (a => 157, b => 226, p => True ), (a => 158, b => 225, p => True ), (a => 159, b => 224, p => True ), (a => 160, b => 223, p => True ), (a => 161, b => 222, p => True ), (a => 162, b => 221, p => True ), (a => 163, b => 220, p => True ), (a => 188, b => 195, p => True ), (a => 189, b => 194, p => True ), (a => 190, b => 193, p => True ), (a => 191, b => 192, p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 40 , b => 48 , p => False), (a => 12 , b => 20 , p => False), (a => 44 , b => 52 , p => False), (a => 10 , b => 18 , p => False), (a => 42 , b => 50 , p => False), (a => 14 , b => 22 , p => False), (a => 46 , b => 54 , p => False), (a => 9  , b => 17 , p => False), (a => 41 , b => 49 , p => False), (a => 13 , b => 21 , p => False), (a => 45 , b => 53 , p => False), (a => 11 , b => 19 , p => False), (a => 43 , b => 51 , p => False), (a => 15 , b => 23 , p => False), (a => 47 , b => 55 , p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 78 , b => 80 , p => False), (a => 82 , b => 84 , p => False), (a => 86 , b => 88 , p => False), (a => 90 , b => 92 , p => False), (a => 98 , b => 100, p => False), (a => 102, b => 104, p => False), (a => 106, b => 108, p => False), (a => 110, b => 112, p => False), (a => 114, b => 116, p => False), (a => 118, b => 120, p => False), (a => 122, b => 124, p => False), (a => 130, b => 132, p => False), (a => 134, b => 136, p => False), (a => 138, b => 140, p => False), (a => 142, b => 144, p => False), (a => 146, b => 148, p => False), (a => 150, b => 152, p => False), (a => 154, b => 156, p => False), (a => 162, b => 164, p => False), (a => 166, b => 168, p => False), (a => 170, b => 172, p => False), (a => 174, b => 176, p => False), (a => 178, b => 180, p => False), (a => 182, b => 184, p => False), (a => 186, b => 188, p => False), (a => 194, b => 196, p => False), (a => 198, b => 200, p => False), (a => 202, b => 204, p => False), (a => 206, b => 208, p => False), (a => 210, b => 212, p => False), (a => 214, b => 216, p => False), (a => 218, b => 220, p => False), (a => 226, b => 228, p => False), (a => 230, b => 232, p => False), (a => 234, b => 236, p => False), (a => 238, b => 240, p => False), (a => 242, b => 244, p => False), (a => 246, b => 248, p => False), (a => 250, b => 252, p => False), (a => 258, b => 260, p => False), (a => 262, b => 264, p => False), (a => 266, b => 268, p => False), (a => 270, b => 272, p => False), (a => 274, b => 276, p => False), (a => 278, b => 280, p => False), (a => 282, b => 284, p => False), (a => 290, b => 292, p => False), (a => 294, b => 296, p => False), (a => 298, b => 300, p => False), (a => 302, b => 304, p => False), (a => 306, b => 308, p => False), (a => 310, b => 312, p => False), (a => 314, b => 316, p => False), (a => 322, b => 324, p => False), (a => 326, b => 328, p => False), (a => 330, b => 332, p => False), (a => 334, b => 336, p => False), (a => 338, b => 340, p => False), (a => 342, b => 344, p => False), (a => 346, b => 348, p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 79 , b => 81 , p => False), (a => 83 , b => 85 , p => False), (a => 87 , b => 89 , p => False), (a => 91 , b => 93 , p => False), (a => 99 , b => 101, p => False), (a => 103, b => 105, p => False), (a => 107, b => 109, p => False), (a => 111, b => 113, p => False), (a => 115, b => 117, p => False), (a => 119, b => 121, p => False), (a => 123, b => 125, p => False), (a => 131, b => 133, p => False), (a => 135, b => 137, p => False), (a => 139, b => 141, p => False), (a => 143, b => 145, p => False), (a => 147, b => 149, p => False), (a => 151, b => 153, p => False), (a => 155, b => 157, p => False), (a => 163, b => 165, p => False), (a => 167, b => 169, p => False), (a => 171, b => 173, p => False), (a => 175, b => 177, p => False), (a => 179, b => 181, p => False), (a => 183, b => 185, p => False), (a => 187, b => 189, p => False), (a => 195, b => 197, p => False), (a => 199, b => 201, p => False), (a => 203, b => 205, p => False), (a => 207, b => 209, p => False), (a => 211, b => 213, p => False), (a => 215, b => 217, p => False), (a => 219, b => 221, p => False), (a => 227, b => 229, p => False), (a => 231, b => 233, p => False), (a => 235, b => 237, p => False), (a => 239, b => 241, p => False), (a => 243, b => 245, p => False), (a => 247, b => 249, p => False), (a => 251, b => 253, p => False), (a => 259, b => 261, p => False), (a => 263, b => 265, p => False), (a => 267, b => 269, p => False), (a => 271, b => 273, p => False), (a => 275, b => 277, p => False), (a => 279, b => 281, p => False), (a => 283, b => 285, p => False), (a => 291, b => 293, p => False), (a => 295, b => 297, p => False), (a => 299, b => 301, p => False), (a => 303, b => 305, p => False), (a => 307, b => 309, p => False), (a => 311, b => 313, p => False), (a => 315, b => 317, p => False), (a => 323, b => 325, p => False), (a => 327, b => 329, p => False), (a => 331, b => 333, p => False), (a => 335, b => 337, p => False), (a => 339, b => 341, p => False), (a => 343, b => 345, p => False), (a => 347, b => 349, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 321, p => True ), (a => 3  , b => 320, p => True ), (a => 4  , b => 319, p => True ), (a => 5  , b => 318, p => True ), (a => 6  , b => 289, p => True ), (a => 7  , b => 288, p => True ), (a => 24 , b => 287, p => True ), (a => 25 , b => 286, p => True ), (a => 26 , b => 257, p => True ), (a => 27 , b => 256, p => True ), (a => 28 , b => 255, p => True ), (a => 29 , b => 254, p => True ), (a => 30 , b => 225, p => True ), (a => 31 , b => 224, p => True ), (a => 32 , b => 223, p => True ), (a => 33 , b => 222, p => True ), (a => 34 , b => 193, p => True ), (a => 35 , b => 192, p => True ), (a => 36 , b => 191, p => True ), (a => 37 , b => 190, p => True ), (a => 38 , b => 161, p => True ), (a => 39 , b => 160, p => True ), (a => 56 , b => 159, p => True ), (a => 57 , b => 158, p => True ), (a => 58 , b => 129, p => True ), (a => 59 , b => 128, p => True ), (a => 60 , b => 127, p => True ), (a => 61 , b => 126, p => True ), (a => 62 , b => 97 , p => True ), (a => 63 , b => 96 , p => True ), (a => 64 , b => 95 , p => True ), (a => 65 , b => 94 , p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 36 , b => 40 , p => False), (a => 44 , b => 48 , p => False), (a => 52 , b => 56 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 38 , b => 42 , p => False), (a => 46 , b => 50 , p => False), (a => 54 , b => 58 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 37 , b => 41 , p => False), (a => 45 , b => 49 , p => False), (a => 53 , b => 57 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 39 , b => 43 , p => False), (a => 47 , b => 51 , p => False), (a => 55 , b => 59 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 79 , b => 80 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 87 , b => 88 , p => False), (a => 89 , b => 90 , p => False), (a => 91 , b => 92 , p => False), (a => 93 , b => 94 , p => False), (a => 97 , b => 98 , p => False), (a => 99 , b => 100, p => False), (a => 101, b => 102, p => False), (a => 103, b => 104, p => False), (a => 105, b => 106, p => False), (a => 107, b => 108, p => False), (a => 109, b => 110, p => False), (a => 111, b => 112, p => False), (a => 113, b => 114, p => False), (a => 115, b => 116, p => False), (a => 117, b => 118, p => False), (a => 119, b => 120, p => False), (a => 121, b => 122, p => False), (a => 123, b => 124, p => False), (a => 125, b => 126, p => False), (a => 129, b => 130, p => False), (a => 131, b => 132, p => False), (a => 133, b => 134, p => False), (a => 135, b => 136, p => False), (a => 137, b => 138, p => False), (a => 139, b => 140, p => False), (a => 141, b => 142, p => False), (a => 143, b => 144, p => False), (a => 145, b => 146, p => False), (a => 147, b => 148, p => False), (a => 149, b => 150, p => False), (a => 151, b => 152, p => False), (a => 153, b => 154, p => False), (a => 155, b => 156, p => False), (a => 157, b => 158, p => False), (a => 161, b => 162, p => False), (a => 163, b => 164, p => False), (a => 165, b => 166, p => False), (a => 167, b => 168, p => False), (a => 169, b => 170, p => False), (a => 171, b => 172, p => False), (a => 173, b => 174, p => False), (a => 175, b => 176, p => False), (a => 177, b => 178, p => False), (a => 179, b => 180, p => False), (a => 181, b => 182, p => False), (a => 183, b => 184, p => False), (a => 185, b => 186, p => False), (a => 187, b => 188, p => False), (a => 189, b => 190, p => False), (a => 193, b => 194, p => False), (a => 195, b => 196, p => False), (a => 197, b => 198, p => False), (a => 199, b => 200, p => False), (a => 201, b => 202, p => False), (a => 203, b => 204, p => False), (a => 205, b => 206, p => False), (a => 207, b => 208, p => False), (a => 209, b => 210, p => False), (a => 211, b => 212, p => False), (a => 213, b => 214, p => False), (a => 215, b => 216, p => False), (a => 217, b => 218, p => False), (a => 219, b => 220, p => False), (a => 221, b => 222, p => False), (a => 225, b => 226, p => False), (a => 227, b => 228, p => False), (a => 229, b => 230, p => False), (a => 231, b => 232, p => False), (a => 233, b => 234, p => False), (a => 235, b => 236, p => False), (a => 237, b => 238, p => False), (a => 239, b => 240, p => False), (a => 241, b => 242, p => False), (a => 243, b => 244, p => False), (a => 245, b => 246, p => False), (a => 247, b => 248, p => False), (a => 249, b => 250, p => False), (a => 251, b => 252, p => False), (a => 253, b => 254, p => False), (a => 257, b => 258, p => False), (a => 259, b => 260, p => False), (a => 261, b => 262, p => False), (a => 263, b => 264, p => False), (a => 265, b => 266, p => False), (a => 267, b => 268, p => False), (a => 269, b => 270, p => False), (a => 271, b => 272, p => False), (a => 273, b => 274, p => False), (a => 275, b => 276, p => False), (a => 277, b => 278, p => False), (a => 279, b => 280, p => False), (a => 281, b => 282, p => False), (a => 283, b => 284, p => False), (a => 285, b => 286, p => False), (a => 289, b => 290, p => False), (a => 291, b => 292, p => False), (a => 293, b => 294, p => False), (a => 295, b => 296, p => False), (a => 297, b => 298, p => False), (a => 299, b => 300, p => False), (a => 301, b => 302, p => False), (a => 303, b => 304, p => False), (a => 305, b => 306, p => False), (a => 307, b => 308, p => False), (a => 309, b => 310, p => False), (a => 311, b => 312, p => False), (a => 313, b => 314, p => False), (a => 315, b => 316, p => False), (a => 317, b => 318, p => False), (a => 321, b => 322, p => False), (a => 323, b => 324, p => False), (a => 325, b => 326, p => False), (a => 327, b => 328, p => False), (a => 329, b => 330, p => False), (a => 331, b => 332, p => False), (a => 333, b => 334, p => False), (a => 335, b => 336, p => False), (a => 337, b => 338, p => False), (a => 339, b => 340, p => False), (a => 341, b => 342, p => False), (a => 343, b => 344, p => False), (a => 345, b => 346, p => False), (a => 347, b => 348, p => False), (a => 349, b => 350, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 320, p => True ), (a => 2  , b => 319, p => True ), (a => 3  , b => 288, p => True ), (a => 28 , b => 287, p => True ), (a => 29 , b => 256, p => True ), (a => 30 , b => 255, p => True ), (a => 31 , b => 224, p => True ), (a => 32 , b => 223, p => True ), (a => 33 , b => 192, p => True ), (a => 34 , b => 191, p => True ), (a => 35 , b => 160, p => True ), (a => 60 , b => 159, p => True ), (a => 61 , b => 128, p => True ), (a => 62 , b => 127, p => True ), (a => 63 , b => 96 , p => True ), (a => 64 , b => 95 , p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 46 , b => 48 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 47 , b => 49 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 80 , b => 112, p => False), (a => 144, b => 176, p => False), (a => 208, b => 240, p => False), (a => 272, b => 304, p => False), (a => 72 , b => 104, p => False), (a => 136, b => 168, p => False), (a => 200, b => 232, p => False), (a => 264, b => 296, p => False), (a => 88 , b => 120, p => False), (a => 152, b => 184, p => False), (a => 216, b => 248, p => False), (a => 280, b => 312, p => False), (a => 68 , b => 100, p => False), (a => 132, b => 164, p => False), (a => 196, b => 228, p => False), (a => 260, b => 292, p => False), (a => 84 , b => 116, p => False), (a => 148, b => 180, p => False), (a => 212, b => 244, p => False), (a => 276, b => 308, p => False), (a => 76 , b => 108, p => False), (a => 140, b => 172, p => False), (a => 204, b => 236, p => False), (a => 268, b => 300, p => False), (a => 92 , b => 124, p => False), (a => 156, b => 188, p => False), (a => 220, b => 252, p => False), (a => 284, b => 316, p => False), (a => 66 , b => 98 , p => False), (a => 130, b => 162, p => False), (a => 194, b => 226, p => False), (a => 258, b => 290, p => False), (a => 82 , b => 114, p => False), (a => 146, b => 178, p => False), (a => 210, b => 242, p => False), (a => 274, b => 306, p => False), (a => 74 , b => 106, p => False), (a => 138, b => 170, p => False), (a => 202, b => 234, p => False), (a => 266, b => 298, p => False), (a => 90 , b => 122, p => False), (a => 154, b => 186, p => False), (a => 218, b => 250, p => False), (a => 282, b => 314, p => False), (a => 70 , b => 102, p => False), (a => 134, b => 166, p => False), (a => 198, b => 230, p => False), (a => 262, b => 294, p => False), (a => 86 , b => 118, p => False), (a => 150, b => 182, p => False), (a => 214, b => 246, p => False), (a => 278, b => 310, p => False), (a => 78 , b => 110, p => False), (a => 142, b => 174, p => False), (a => 206, b => 238, p => False), (a => 270, b => 302, p => False), (a => 94 , b => 126, p => False), (a => 158, b => 190, p => False), (a => 222, b => 254, p => False), (a => 286, b => 318, p => False), (a => 65 , b => 97 , p => False), (a => 129, b => 161, p => False), (a => 193, b => 225, p => False), (a => 257, b => 289, p => False), (a => 81 , b => 113, p => False), (a => 145, b => 177, p => False), (a => 209, b => 241, p => False), (a => 273, b => 305, p => False), (a => 73 , b => 105, p => False), (a => 137, b => 169, p => False), (a => 201, b => 233, p => False), (a => 265, b => 297, p => False), (a => 89 , b => 121, p => False), (a => 153, b => 185, p => False), (a => 217, b => 249, p => False), (a => 281, b => 313, p => False), (a => 69 , b => 101, p => False), (a => 133, b => 165, p => False), (a => 197, b => 229, p => False), (a => 261, b => 293, p => False), (a => 85 , b => 117, p => False), (a => 149, b => 181, p => False), (a => 213, b => 245, p => False), (a => 277, b => 309, p => False), (a => 77 , b => 109, p => False), (a => 141, b => 173, p => False), (a => 205, b => 237, p => False), (a => 269, b => 301, p => False), (a => 93 , b => 125, p => False), (a => 157, b => 189, p => False), (a => 221, b => 253, p => False), (a => 285, b => 317, p => False), (a => 67 , b => 99 , p => False), (a => 131, b => 163, p => False), (a => 195, b => 227, p => False), (a => 259, b => 291, p => False), (a => 83 , b => 115, p => False), (a => 147, b => 179, p => False), (a => 211, b => 243, p => False), (a => 275, b => 307, p => False), (a => 75 , b => 107, p => False), (a => 139, b => 171, p => False), (a => 203, b => 235, p => False), (a => 267, b => 299, p => False), (a => 91 , b => 123, p => False), (a => 155, b => 187, p => False), (a => 219, b => 251, p => False), (a => 283, b => 315, p => False), (a => 71 , b => 103, p => False), (a => 135, b => 167, p => False), (a => 199, b => 231, p => False), (a => 263, b => 295, p => False), (a => 87 , b => 119, p => False), (a => 151, b => 183, p => False), (a => 215, b => 247, p => False), (a => 279, b => 311, p => False), (a => 79 , b => 111, p => False), (a => 143, b => 175, p => False), (a => 207, b => 239, p => False), (a => 271, b => 303, p => False), (a => 328, b => 336, p => False), (a => 332, b => 340, p => False), (a => 330, b => 338, p => False), (a => 334, b => 342, p => False), (a => 329, b => 337, p => False), (a => 333, b => 341, p => False), (a => 331, b => 339, p => False), (a => 335, b => 343, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 30 , b => 349, p => True ), (a => 31 , b => 348, p => True ), (a => 32 , b => 347, p => True ), (a => 33 , b => 346, p => True ), (a => 62 , b => 345, p => True ), (a => 63 , b => 344, p => True ), (a => 64 , b => 327, p => True ), (a => 95 , b => 326, p => True ), (a => 96 , b => 325, p => True ), (a => 127, b => 324, p => True ), (a => 128, b => 323, p => True ), (a => 159, b => 322, p => True ), (a => 160, b => 321, p => True ), (a => 191, b => 320, p => True ), (a => 192, b => 319, p => True ), (a => 223, b => 288, p => True ), (a => 224, b => 287, p => True ), (a => 255, b => 256, p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 47 , b => 48 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 80 , b => 96 , p => False), (a => 144, b => 160, p => False), (a => 208, b => 224, p => False), (a => 272, b => 288, p => False), (a => 88 , b => 104, p => False), (a => 152, b => 168, p => False), (a => 216, b => 232, p => False), (a => 280, b => 296, p => False), (a => 84 , b => 100, p => False), (a => 148, b => 164, p => False), (a => 212, b => 228, p => False), (a => 276, b => 292, p => False), (a => 92 , b => 108, p => False), (a => 156, b => 172, p => False), (a => 220, b => 236, p => False), (a => 284, b => 300, p => False), (a => 82 , b => 98 , p => False), (a => 146, b => 162, p => False), (a => 210, b => 226, p => False), (a => 274, b => 290, p => False), (a => 90 , b => 106, p => False), (a => 154, b => 170, p => False), (a => 218, b => 234, p => False), (a => 282, b => 298, p => False), (a => 86 , b => 102, p => False), (a => 150, b => 166, p => False), (a => 214, b => 230, p => False), (a => 278, b => 294, p => False), (a => 94 , b => 110, p => False), (a => 158, b => 174, p => False), (a => 222, b => 238, p => False), (a => 286, b => 302, p => False), (a => 81 , b => 97 , p => False), (a => 145, b => 161, p => False), (a => 209, b => 225, p => False), (a => 273, b => 289, p => False), (a => 89 , b => 105, p => False), (a => 153, b => 169, p => False), (a => 217, b => 233, p => False), (a => 281, b => 297, p => False), (a => 85 , b => 101, p => False), (a => 149, b => 165, p => False), (a => 213, b => 229, p => False), (a => 277, b => 293, p => False), (a => 93 , b => 109, p => False), (a => 157, b => 173, p => False), (a => 221, b => 237, p => False), (a => 285, b => 301, p => False), (a => 83 , b => 99 , p => False), (a => 147, b => 163, p => False), (a => 211, b => 227, p => False), (a => 275, b => 291, p => False), (a => 91 , b => 107, p => False), (a => 155, b => 171, p => False), (a => 219, b => 235, p => False), (a => 283, b => 299, p => False), (a => 87 , b => 103, p => False), (a => 151, b => 167, p => False), (a => 215, b => 231, p => False), (a => 279, b => 295, p => False), (a => 95 , b => 111, p => False), (a => 159, b => 175, p => False), (a => 223, b => 239, p => False), (a => 287, b => 303, p => False), (a => 324, b => 328, p => False), (a => 332, b => 336, p => False), (a => 340, b => 344, p => False), (a => 326, b => 330, p => False), (a => 334, b => 338, p => False), (a => 342, b => 346, p => False), (a => 325, b => 329, p => False), (a => 333, b => 337, p => False), (a => 341, b => 345, p => False), (a => 327, b => 331, p => False), (a => 335, b => 339, p => False), (a => 343, b => 347, p => False), (a => 0  , b => 351, p => True ), (a => 31 , b => 350, p => True ), (a => 32 , b => 349, p => True ), (a => 63 , b => 348, p => True ), (a => 64 , b => 323, p => True ), (a => 65 , b => 322, p => True ), (a => 66 , b => 321, p => True ), (a => 67 , b => 320, p => True ), (a => 68 , b => 319, p => True ), (a => 69 , b => 318, p => True ), (a => 70 , b => 317, p => True ), (a => 71 , b => 316, p => True ), (a => 72 , b => 315, p => True ), (a => 73 , b => 314, p => True ), (a => 74 , b => 313, p => True ), (a => 75 , b => 312, p => True ), (a => 76 , b => 311, p => True ), (a => 77 , b => 310, p => True ), (a => 78 , b => 309, p => True ), (a => 79 , b => 308, p => True ), (a => 112, b => 307, p => True ), (a => 113, b => 306, p => True ), (a => 114, b => 305, p => True ), (a => 115, b => 304, p => True ), (a => 116, b => 271, p => True ), (a => 117, b => 270, p => True ), (a => 118, b => 269, p => True ), (a => 119, b => 268, p => True ), (a => 120, b => 267, p => True ), (a => 121, b => 266, p => True ), (a => 122, b => 265, p => True ), (a => 123, b => 264, p => True ), (a => 124, b => 263, p => True ), (a => 125, b => 262, p => True ), (a => 126, b => 261, p => True ), (a => 127, b => 260, p => True ), (a => 128, b => 259, p => True ), (a => 129, b => 258, p => True ), (a => 130, b => 257, p => True ), (a => 131, b => 256, p => True ), (a => 132, b => 255, p => True ), (a => 133, b => 254, p => True ), (a => 134, b => 253, p => True ), (a => 135, b => 252, p => True ), (a => 136, b => 251, p => True ), (a => 137, b => 250, p => True ), (a => 138, b => 249, p => True ), (a => 139, b => 248, p => True ), (a => 140, b => 247, p => True ), (a => 141, b => 246, p => True ), (a => 142, b => 245, p => True ), (a => 143, b => 244, p => True ), (a => 176, b => 243, p => True ), (a => 177, b => 242, p => True ), (a => 178, b => 241, p => True ), (a => 179, b => 240, p => True ), (a => 180, b => 207, p => True ), (a => 181, b => 206, p => True ), (a => 182, b => 205, p => True ), (a => 183, b => 204, p => True ), (a => 184, b => 203, p => True ), (a => 185, b => 202, p => True ), (a => 186, b => 201, p => True ), (a => 187, b => 200, p => True ), (a => 188, b => 199, p => True ), (a => 189, b => 198, p => True ), (a => 190, b => 197, p => True ), (a => 191, b => 196, p => True ), (a => 192, b => 195, p => True ), (a => 193, b => 194, p => True )),
                    ((a => 16 , b => 48 , p => False), (a => 8  , b => 40 , p => False), (a => 24 , b => 56 , p => False), (a => 4  , b => 36 , p => False), (a => 20 , b => 52 , p => False), (a => 12 , b => 44 , p => False), (a => 28 , b => 60 , p => False), (a => 2  , b => 34 , p => False), (a => 18 , b => 50 , p => False), (a => 10 , b => 42 , p => False), (a => 26 , b => 58 , p => False), (a => 6  , b => 38 , p => False), (a => 22 , b => 54 , p => False), (a => 14 , b => 46 , p => False), (a => 30 , b => 62 , p => False), (a => 1  , b => 33 , p => False), (a => 17 , b => 49 , p => False), (a => 9  , b => 41 , p => False), (a => 25 , b => 57 , p => False), (a => 5  , b => 37 , p => False), (a => 21 , b => 53 , p => False), (a => 13 , b => 45 , p => False), (a => 29 , b => 61 , p => False), (a => 3  , b => 35 , p => False), (a => 19 , b => 51 , p => False), (a => 11 , b => 43 , p => False), (a => 27 , b => 59 , p => False), (a => 7  , b => 39 , p => False), (a => 23 , b => 55 , p => False), (a => 15 , b => 47 , p => False), (a => 72 , b => 80 , p => False), (a => 88 , b => 96 , p => False), (a => 104, b => 112, p => False), (a => 136, b => 144, p => False), (a => 152, b => 160, p => False), (a => 168, b => 176, p => False), (a => 200, b => 208, p => False), (a => 216, b => 224, p => False), (a => 232, b => 240, p => False), (a => 264, b => 272, p => False), (a => 280, b => 288, p => False), (a => 296, b => 304, p => False), (a => 76 , b => 84 , p => False), (a => 92 , b => 100, p => False), (a => 108, b => 116, p => False), (a => 140, b => 148, p => False), (a => 156, b => 164, p => False), (a => 172, b => 180, p => False), (a => 204, b => 212, p => False), (a => 220, b => 228, p => False), (a => 236, b => 244, p => False), (a => 268, b => 276, p => False), (a => 284, b => 292, p => False), (a => 300, b => 308, p => False), (a => 74 , b => 82 , p => False), (a => 90 , b => 98 , p => False), (a => 106, b => 114, p => False), (a => 138, b => 146, p => False), (a => 154, b => 162, p => False), (a => 170, b => 178, p => False), (a => 202, b => 210, p => False), (a => 218, b => 226, p => False), (a => 234, b => 242, p => False), (a => 266, b => 274, p => False), (a => 282, b => 290, p => False), (a => 298, b => 306, p => False), (a => 78 , b => 86 , p => False), (a => 94 , b => 102, p => False), (a => 110, b => 118, p => False), (a => 142, b => 150, p => False), (a => 158, b => 166, p => False), (a => 174, b => 182, p => False), (a => 206, b => 214, p => False), (a => 222, b => 230, p => False), (a => 238, b => 246, p => False), (a => 270, b => 278, p => False), (a => 286, b => 294, p => False), (a => 302, b => 310, p => False), (a => 73 , b => 81 , p => False), (a => 89 , b => 97 , p => False), (a => 105, b => 113, p => False), (a => 137, b => 145, p => False), (a => 153, b => 161, p => False), (a => 169, b => 177, p => False), (a => 201, b => 209, p => False), (a => 217, b => 225, p => False), (a => 233, b => 241, p => False), (a => 265, b => 273, p => False), (a => 281, b => 289, p => False), (a => 297, b => 305, p => False), (a => 77 , b => 85 , p => False), (a => 93 , b => 101, p => False), (a => 109, b => 117, p => False), (a => 141, b => 149, p => False), (a => 157, b => 165, p => False), (a => 173, b => 181, p => False), (a => 205, b => 213, p => False), (a => 221, b => 229, p => False), (a => 237, b => 245, p => False), (a => 269, b => 277, p => False), (a => 285, b => 293, p => False), (a => 301, b => 309, p => False), (a => 75 , b => 83 , p => False), (a => 91 , b => 99 , p => False), (a => 107, b => 115, p => False), (a => 139, b => 147, p => False), (a => 155, b => 163, p => False), (a => 171, b => 179, p => False), (a => 203, b => 211, p => False), (a => 219, b => 227, p => False), (a => 235, b => 243, p => False), (a => 267, b => 275, p => False), (a => 283, b => 291, p => False), (a => 299, b => 307, p => False), (a => 79 , b => 87 , p => False), (a => 95 , b => 103, p => False), (a => 111, b => 119, p => False), (a => 143, b => 151, p => False), (a => 159, b => 167, p => False), (a => 175, b => 183, p => False), (a => 207, b => 215, p => False), (a => 223, b => 231, p => False), (a => 239, b => 247, p => False), (a => 271, b => 279, p => False), (a => 287, b => 295, p => False), (a => 303, b => 311, p => False), (a => 322, b => 324, p => False), (a => 326, b => 328, p => False), (a => 330, b => 332, p => False), (a => 334, b => 336, p => False), (a => 338, b => 340, p => False), (a => 342, b => 344, p => False), (a => 346, b => 348, p => False), (a => 323, b => 325, p => False), (a => 327, b => 329, p => False), (a => 331, b => 333, p => False), (a => 335, b => 337, p => False), (a => 339, b => 341, p => False), (a => 343, b => 345, p => False), (a => 347, b => 349, p => False), (a => 0  , b => 351, p => True ), (a => 31 , b => 350, p => True ), (a => 32 , b => 321, p => True ), (a => 63 , b => 320, p => True ), (a => 64 , b => 319, p => True ), (a => 65 , b => 318, p => True ), (a => 66 , b => 317, p => True ), (a => 67 , b => 316, p => True ), (a => 68 , b => 315, p => True ), (a => 69 , b => 314, p => True ), (a => 70 , b => 313, p => True ), (a => 71 , b => 312, p => True ), (a => 120, b => 263, p => True ), (a => 121, b => 262, p => True ), (a => 122, b => 261, p => True ), (a => 123, b => 260, p => True ), (a => 124, b => 259, p => True ), (a => 125, b => 258, p => True ), (a => 126, b => 257, p => True ), (a => 127, b => 256, p => True ), (a => 128, b => 255, p => True ), (a => 129, b => 254, p => True ), (a => 130, b => 253, p => True ), (a => 131, b => 252, p => True ), (a => 132, b => 251, p => True ), (a => 133, b => 250, p => True ), (a => 134, b => 249, p => True ), (a => 135, b => 248, p => True ), (a => 184, b => 199, p => True ), (a => 185, b => 198, p => True ), (a => 186, b => 197, p => True ), (a => 187, b => 196, p => True ), (a => 188, b => 195, p => True ), (a => 189, b => 194, p => True ), (a => 190, b => 193, p => True ), (a => 191, b => 192, p => True )),
                    ((a => 16 , b => 32 , p => False), (a => 24 , b => 40 , p => False), (a => 20 , b => 36 , p => False), (a => 28 , b => 44 , p => False), (a => 18 , b => 34 , p => False), (a => 26 , b => 42 , p => False), (a => 22 , b => 38 , p => False), (a => 30 , b => 46 , p => False), (a => 17 , b => 33 , p => False), (a => 25 , b => 41 , p => False), (a => 21 , b => 37 , p => False), (a => 29 , b => 45 , p => False), (a => 19 , b => 35 , p => False), (a => 27 , b => 43 , p => False), (a => 23 , b => 39 , p => False), (a => 31 , b => 47 , p => False), (a => 68 , b => 72 , p => False), (a => 76 , b => 80 , p => False), (a => 84 , b => 88 , p => False), (a => 92 , b => 96 , p => False), (a => 100, b => 104, p => False), (a => 108, b => 112, p => False), (a => 116, b => 120, p => False), (a => 132, b => 136, p => False), (a => 140, b => 144, p => False), (a => 148, b => 152, p => False), (a => 156, b => 160, p => False), (a => 164, b => 168, p => False), (a => 172, b => 176, p => False), (a => 180, b => 184, p => False), (a => 196, b => 200, p => False), (a => 204, b => 208, p => False), (a => 212, b => 216, p => False), (a => 220, b => 224, p => False), (a => 228, b => 232, p => False), (a => 236, b => 240, p => False), (a => 244, b => 248, p => False), (a => 260, b => 264, p => False), (a => 268, b => 272, p => False), (a => 276, b => 280, p => False), (a => 284, b => 288, p => False), (a => 292, b => 296, p => False), (a => 300, b => 304, p => False), (a => 308, b => 312, p => False), (a => 70 , b => 74 , p => False), (a => 78 , b => 82 , p => False), (a => 86 , b => 90 , p => False), (a => 94 , b => 98 , p => False), (a => 102, b => 106, p => False), (a => 110, b => 114, p => False), (a => 118, b => 122, p => False), (a => 134, b => 138, p => False), (a => 142, b => 146, p => False), (a => 150, b => 154, p => False), (a => 158, b => 162, p => False), (a => 166, b => 170, p => False), (a => 174, b => 178, p => False), (a => 182, b => 186, p => False), (a => 198, b => 202, p => False), (a => 206, b => 210, p => False), (a => 214, b => 218, p => False), (a => 222, b => 226, p => False), (a => 230, b => 234, p => False), (a => 238, b => 242, p => False), (a => 246, b => 250, p => False), (a => 262, b => 266, p => False), (a => 270, b => 274, p => False), (a => 278, b => 282, p => False), (a => 286, b => 290, p => False), (a => 294, b => 298, p => False), (a => 302, b => 306, p => False), (a => 310, b => 314, p => False), (a => 69 , b => 73 , p => False), (a => 77 , b => 81 , p => False), (a => 85 , b => 89 , p => False), (a => 93 , b => 97 , p => False), (a => 101, b => 105, p => False), (a => 109, b => 113, p => False), (a => 117, b => 121, p => False), (a => 133, b => 137, p => False), (a => 141, b => 145, p => False), (a => 149, b => 153, p => False), (a => 157, b => 161, p => False), (a => 165, b => 169, p => False), (a => 173, b => 177, p => False), (a => 181, b => 185, p => False), (a => 197, b => 201, p => False), (a => 205, b => 209, p => False), (a => 213, b => 217, p => False), (a => 221, b => 225, p => False), (a => 229, b => 233, p => False), (a => 237, b => 241, p => False), (a => 245, b => 249, p => False), (a => 261, b => 265, p => False), (a => 269, b => 273, p => False), (a => 277, b => 281, p => False), (a => 285, b => 289, p => False), (a => 293, b => 297, p => False), (a => 301, b => 305, p => False), (a => 309, b => 313, p => False), (a => 71 , b => 75 , p => False), (a => 79 , b => 83 , p => False), (a => 87 , b => 91 , p => False), (a => 95 , b => 99 , p => False), (a => 103, b => 107, p => False), (a => 111, b => 115, p => False), (a => 119, b => 123, p => False), (a => 135, b => 139, p => False), (a => 143, b => 147, p => False), (a => 151, b => 155, p => False), (a => 159, b => 163, p => False), (a => 167, b => 171, p => False), (a => 175, b => 179, p => False), (a => 183, b => 187, p => False), (a => 199, b => 203, p => False), (a => 207, b => 211, p => False), (a => 215, b => 219, p => False), (a => 223, b => 227, p => False), (a => 231, b => 235, p => False), (a => 239, b => 243, p => False), (a => 247, b => 251, p => False), (a => 263, b => 267, p => False), (a => 271, b => 275, p => False), (a => 279, b => 283, p => False), (a => 287, b => 291, p => False), (a => 295, b => 299, p => False), (a => 303, b => 307, p => False), (a => 311, b => 315, p => False), (a => 321, b => 322, p => False), (a => 323, b => 324, p => False), (a => 325, b => 326, p => False), (a => 327, b => 328, p => False), (a => 329, b => 330, p => False), (a => 331, b => 332, p => False), (a => 333, b => 334, p => False), (a => 335, b => 336, p => False), (a => 337, b => 338, p => False), (a => 339, b => 340, p => False), (a => 341, b => 342, p => False), (a => 343, b => 344, p => False), (a => 345, b => 346, p => False), (a => 347, b => 348, p => False), (a => 349, b => 350, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 320, p => True ), (a => 2  , b => 319, p => True ), (a => 3  , b => 318, p => True ), (a => 4  , b => 317, p => True ), (a => 5  , b => 316, p => True ), (a => 6  , b => 259, p => True ), (a => 7  , b => 258, p => True ), (a => 8  , b => 257, p => True ), (a => 9  , b => 256, p => True ), (a => 10 , b => 255, p => True ), (a => 11 , b => 254, p => True ), (a => 12 , b => 253, p => True ), (a => 13 , b => 252, p => True ), (a => 14 , b => 195, p => True ), (a => 15 , b => 194, p => True ), (a => 48 , b => 193, p => True ), (a => 49 , b => 192, p => True ), (a => 50 , b => 191, p => True ), (a => 51 , b => 190, p => True ), (a => 52 , b => 189, p => True ), (a => 53 , b => 188, p => True ), (a => 54 , b => 131, p => True ), (a => 55 , b => 130, p => True ), (a => 56 , b => 129, p => True ), (a => 57 , b => 128, p => True ), (a => 58 , b => 127, p => True ), (a => 59 , b => 126, p => True ), (a => 60 , b => 125, p => True ), (a => 61 , b => 124, p => True ), (a => 62 , b => 67 , p => True ), (a => 63 , b => 66 , p => True ), (a => 64 , b => 65 , p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 24 , b => 32 , p => False), (a => 40 , b => 48 , p => False), (a => 12 , b => 20 , p => False), (a => 28 , b => 36 , p => False), (a => 44 , b => 52 , p => False), (a => 10 , b => 18 , p => False), (a => 26 , b => 34 , p => False), (a => 42 , b => 50 , p => False), (a => 14 , b => 22 , p => False), (a => 30 , b => 38 , p => False), (a => 46 , b => 54 , p => False), (a => 9  , b => 17 , p => False), (a => 25 , b => 33 , p => False), (a => 41 , b => 49 , p => False), (a => 13 , b => 21 , p => False), (a => 29 , b => 37 , p => False), (a => 45 , b => 53 , p => False), (a => 11 , b => 19 , p => False), (a => 27 , b => 35 , p => False), (a => 43 , b => 51 , p => False), (a => 15 , b => 23 , p => False), (a => 31 , b => 39 , p => False), (a => 47 , b => 55 , p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 78 , b => 80 , p => False), (a => 82 , b => 84 , p => False), (a => 86 , b => 88 , p => False), (a => 90 , b => 92 , p => False), (a => 94 , b => 96 , p => False), (a => 98 , b => 100, p => False), (a => 102, b => 104, p => False), (a => 106, b => 108, p => False), (a => 110, b => 112, p => False), (a => 114, b => 116, p => False), (a => 118, b => 120, p => False), (a => 122, b => 124, p => False), (a => 130, b => 132, p => False), (a => 134, b => 136, p => False), (a => 138, b => 140, p => False), (a => 142, b => 144, p => False), (a => 146, b => 148, p => False), (a => 150, b => 152, p => False), (a => 154, b => 156, p => False), (a => 158, b => 160, p => False), (a => 162, b => 164, p => False), (a => 166, b => 168, p => False), (a => 170, b => 172, p => False), (a => 174, b => 176, p => False), (a => 178, b => 180, p => False), (a => 182, b => 184, p => False), (a => 186, b => 188, p => False), (a => 194, b => 196, p => False), (a => 198, b => 200, p => False), (a => 202, b => 204, p => False), (a => 206, b => 208, p => False), (a => 210, b => 212, p => False), (a => 214, b => 216, p => False), (a => 218, b => 220, p => False), (a => 222, b => 224, p => False), (a => 226, b => 228, p => False), (a => 230, b => 232, p => False), (a => 234, b => 236, p => False), (a => 238, b => 240, p => False), (a => 242, b => 244, p => False), (a => 246, b => 248, p => False), (a => 250, b => 252, p => False), (a => 258, b => 260, p => False), (a => 262, b => 264, p => False), (a => 266, b => 268, p => False), (a => 270, b => 272, p => False), (a => 274, b => 276, p => False), (a => 278, b => 280, p => False), (a => 282, b => 284, p => False), (a => 286, b => 288, p => False), (a => 290, b => 292, p => False), (a => 294, b => 296, p => False), (a => 298, b => 300, p => False), (a => 302, b => 304, p => False), (a => 306, b => 308, p => False), (a => 310, b => 312, p => False), (a => 314, b => 316, p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 79 , b => 81 , p => False), (a => 83 , b => 85 , p => False), (a => 87 , b => 89 , p => False), (a => 91 , b => 93 , p => False), (a => 95 , b => 97 , p => False), (a => 99 , b => 101, p => False), (a => 103, b => 105, p => False), (a => 107, b => 109, p => False), (a => 111, b => 113, p => False), (a => 115, b => 117, p => False), (a => 119, b => 121, p => False), (a => 123, b => 125, p => False), (a => 131, b => 133, p => False), (a => 135, b => 137, p => False), (a => 139, b => 141, p => False), (a => 143, b => 145, p => False), (a => 147, b => 149, p => False), (a => 151, b => 153, p => False), (a => 155, b => 157, p => False), (a => 159, b => 161, p => False), (a => 163, b => 165, p => False), (a => 167, b => 169, p => False), (a => 171, b => 173, p => False), (a => 175, b => 177, p => False), (a => 179, b => 181, p => False), (a => 183, b => 185, p => False), (a => 187, b => 189, p => False), (a => 195, b => 197, p => False), (a => 199, b => 201, p => False), (a => 203, b => 205, p => False), (a => 207, b => 209, p => False), (a => 211, b => 213, p => False), (a => 215, b => 217, p => False), (a => 219, b => 221, p => False), (a => 223, b => 225, p => False), (a => 227, b => 229, p => False), (a => 231, b => 233, p => False), (a => 235, b => 237, p => False), (a => 239, b => 241, p => False), (a => 243, b => 245, p => False), (a => 247, b => 249, p => False), (a => 251, b => 253, p => False), (a => 259, b => 261, p => False), (a => 263, b => 265, p => False), (a => 267, b => 269, p => False), (a => 271, b => 273, p => False), (a => 275, b => 277, p => False), (a => 279, b => 281, p => False), (a => 283, b => 285, p => False), (a => 287, b => 289, p => False), (a => 291, b => 293, p => False), (a => 295, b => 297, p => False), (a => 299, b => 301, p => False), (a => 303, b => 305, p => False), (a => 307, b => 309, p => False), (a => 311, b => 313, p => False), (a => 315, b => 317, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 56 , b => 343, p => True ), (a => 57 , b => 342, p => True ), (a => 58 , b => 341, p => True ), (a => 59 , b => 340, p => True ), (a => 60 , b => 339, p => True ), (a => 61 , b => 338, p => True ), (a => 62 , b => 337, p => True ), (a => 63 , b => 336, p => True ), (a => 64 , b => 335, p => True ), (a => 65 , b => 334, p => True ), (a => 126, b => 333, p => True ), (a => 127, b => 332, p => True ), (a => 128, b => 331, p => True ), (a => 129, b => 330, p => True ), (a => 190, b => 329, p => True ), (a => 191, b => 328, p => True ), (a => 192, b => 327, p => True ), (a => 193, b => 326, p => True ), (a => 254, b => 325, p => True ), (a => 255, b => 324, p => True ), (a => 256, b => 323, p => True ), (a => 257, b => 322, p => True ), (a => 318, b => 321, p => True ), (a => 319, b => 320, p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 28 , b => 32 , p => False), (a => 36 , b => 40 , p => False), (a => 44 , b => 48 , p => False), (a => 52 , b => 56 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 30 , b => 34 , p => False), (a => 38 , b => 42 , p => False), (a => 46 , b => 50 , p => False), (a => 54 , b => 58 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 29 , b => 33 , p => False), (a => 37 , b => 41 , p => False), (a => 45 , b => 49 , p => False), (a => 53 , b => 57 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 31 , b => 35 , p => False), (a => 39 , b => 43 , p => False), (a => 47 , b => 51 , p => False), (a => 55 , b => 59 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 79 , b => 80 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 87 , b => 88 , p => False), (a => 89 , b => 90 , p => False), (a => 91 , b => 92 , p => False), (a => 93 , b => 94 , p => False), (a => 95 , b => 96 , p => False), (a => 97 , b => 98 , p => False), (a => 99 , b => 100, p => False), (a => 101, b => 102, p => False), (a => 103, b => 104, p => False), (a => 105, b => 106, p => False), (a => 107, b => 108, p => False), (a => 109, b => 110, p => False), (a => 111, b => 112, p => False), (a => 113, b => 114, p => False), (a => 115, b => 116, p => False), (a => 117, b => 118, p => False), (a => 119, b => 120, p => False), (a => 121, b => 122, p => False), (a => 123, b => 124, p => False), (a => 125, b => 126, p => False), (a => 129, b => 130, p => False), (a => 131, b => 132, p => False), (a => 133, b => 134, p => False), (a => 135, b => 136, p => False), (a => 137, b => 138, p => False), (a => 139, b => 140, p => False), (a => 141, b => 142, p => False), (a => 143, b => 144, p => False), (a => 145, b => 146, p => False), (a => 147, b => 148, p => False), (a => 149, b => 150, p => False), (a => 151, b => 152, p => False), (a => 153, b => 154, p => False), (a => 155, b => 156, p => False), (a => 157, b => 158, p => False), (a => 159, b => 160, p => False), (a => 161, b => 162, p => False), (a => 163, b => 164, p => False), (a => 165, b => 166, p => False), (a => 167, b => 168, p => False), (a => 169, b => 170, p => False), (a => 171, b => 172, p => False), (a => 173, b => 174, p => False), (a => 175, b => 176, p => False), (a => 177, b => 178, p => False), (a => 179, b => 180, p => False), (a => 181, b => 182, p => False), (a => 183, b => 184, p => False), (a => 185, b => 186, p => False), (a => 187, b => 188, p => False), (a => 189, b => 190, p => False), (a => 193, b => 194, p => False), (a => 195, b => 196, p => False), (a => 197, b => 198, p => False), (a => 199, b => 200, p => False), (a => 201, b => 202, p => False), (a => 203, b => 204, p => False), (a => 205, b => 206, p => False), (a => 207, b => 208, p => False), (a => 209, b => 210, p => False), (a => 211, b => 212, p => False), (a => 213, b => 214, p => False), (a => 215, b => 216, p => False), (a => 217, b => 218, p => False), (a => 219, b => 220, p => False), (a => 221, b => 222, p => False), (a => 223, b => 224, p => False), (a => 225, b => 226, p => False), (a => 227, b => 228, p => False), (a => 229, b => 230, p => False), (a => 231, b => 232, p => False), (a => 233, b => 234, p => False), (a => 235, b => 236, p => False), (a => 237, b => 238, p => False), (a => 239, b => 240, p => False), (a => 241, b => 242, p => False), (a => 243, b => 244, p => False), (a => 245, b => 246, p => False), (a => 247, b => 248, p => False), (a => 249, b => 250, p => False), (a => 251, b => 252, p => False), (a => 253, b => 254, p => False), (a => 257, b => 258, p => False), (a => 259, b => 260, p => False), (a => 261, b => 262, p => False), (a => 263, b => 264, p => False), (a => 265, b => 266, p => False), (a => 267, b => 268, p => False), (a => 269, b => 270, p => False), (a => 271, b => 272, p => False), (a => 273, b => 274, p => False), (a => 275, b => 276, p => False), (a => 277, b => 278, p => False), (a => 279, b => 280, p => False), (a => 281, b => 282, p => False), (a => 283, b => 284, p => False), (a => 285, b => 286, p => False), (a => 287, b => 288, p => False), (a => 289, b => 290, p => False), (a => 291, b => 292, p => False), (a => 293, b => 294, p => False), (a => 295, b => 296, p => False), (a => 297, b => 298, p => False), (a => 299, b => 300, p => False), (a => 301, b => 302, p => False), (a => 303, b => 304, p => False), (a => 305, b => 306, p => False), (a => 307, b => 308, p => False), (a => 309, b => 310, p => False), (a => 311, b => 312, p => False), (a => 313, b => 314, p => False), (a => 315, b => 316, p => False), (a => 317, b => 318, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 60 , b => 347, p => True ), (a => 61 , b => 346, p => True ), (a => 62 , b => 345, p => True ), (a => 63 , b => 344, p => True ), (a => 64 , b => 343, p => True ), (a => 127, b => 342, p => True ), (a => 128, b => 341, p => True ), (a => 191, b => 340, p => True ), (a => 192, b => 339, p => True ), (a => 255, b => 338, p => True ), (a => 256, b => 337, p => True ), (a => 319, b => 336, p => True ), (a => 320, b => 335, p => True ), (a => 321, b => 334, p => True ), (a => 322, b => 333, p => True ), (a => 323, b => 332, p => True ), (a => 324, b => 331, p => True ), (a => 325, b => 330, p => True ), (a => 326, b => 329, p => True ), (a => 327, b => 328, p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 30 , b => 32 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 46 , b => 48 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 31 , b => 33 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 47 , b => 49 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 160, b => 224, p => False), (a => 144, b => 208, p => False), (a => 272, b => 336, p => False), (a => 176, b => 240, p => False), (a => 136, b => 200, p => False), (a => 264, b => 328, p => False), (a => 168, b => 232, p => False), (a => 152, b => 216, p => False), (a => 280, b => 344, p => False), (a => 184, b => 248, p => False), (a => 132, b => 196, p => False), (a => 260, b => 324, p => False), (a => 164, b => 228, p => False), (a => 148, b => 212, p => False), (a => 276, b => 340, p => False), (a => 180, b => 244, p => False), (a => 140, b => 204, p => False), (a => 268, b => 332, p => False), (a => 172, b => 236, p => False), (a => 156, b => 220, p => False), (a => 284, b => 348, p => False), (a => 188, b => 252, p => False), (a => 130, b => 194, p => False), (a => 258, b => 322, p => False), (a => 162, b => 226, p => False), (a => 146, b => 210, p => False), (a => 274, b => 338, p => False), (a => 178, b => 242, p => False), (a => 138, b => 202, p => False), (a => 266, b => 330, p => False), (a => 170, b => 234, p => False), (a => 154, b => 218, p => False), (a => 282, b => 346, p => False), (a => 186, b => 250, p => False), (a => 134, b => 198, p => False), (a => 262, b => 326, p => False), (a => 166, b => 230, p => False), (a => 150, b => 214, p => False), (a => 278, b => 342, p => False), (a => 182, b => 246, p => False), (a => 142, b => 206, p => False), (a => 270, b => 334, p => False), (a => 174, b => 238, p => False), (a => 158, b => 222, p => False), (a => 286, b => 350, p => False), (a => 190, b => 254, p => False), (a => 129, b => 193, p => False), (a => 257, b => 321, p => False), (a => 161, b => 225, p => False), (a => 145, b => 209, p => False), (a => 273, b => 337, p => False), (a => 177, b => 241, p => False), (a => 137, b => 201, p => False), (a => 265, b => 329, p => False), (a => 169, b => 233, p => False), (a => 153, b => 217, p => False), (a => 281, b => 345, p => False), (a => 185, b => 249, p => False), (a => 133, b => 197, p => False), (a => 261, b => 325, p => False), (a => 165, b => 229, p => False), (a => 149, b => 213, p => False), (a => 277, b => 341, p => False), (a => 181, b => 245, p => False), (a => 141, b => 205, p => False), (a => 269, b => 333, p => False), (a => 173, b => 237, p => False), (a => 157, b => 221, p => False), (a => 285, b => 349, p => False), (a => 189, b => 253, p => False), (a => 131, b => 195, p => False), (a => 259, b => 323, p => False), (a => 163, b => 227, p => False), (a => 147, b => 211, p => False), (a => 275, b => 339, p => False), (a => 179, b => 243, p => False), (a => 139, b => 203, p => False), (a => 267, b => 331, p => False), (a => 171, b => 235, p => False), (a => 155, b => 219, p => False), (a => 283, b => 347, p => False), (a => 187, b => 251, p => False), (a => 135, b => 199, p => False), (a => 263, b => 327, p => False), (a => 167, b => 231, p => False), (a => 151, b => 215, p => False), (a => 279, b => 343, p => False), (a => 183, b => 247, p => False), (a => 143, b => 207, p => False), (a => 271, b => 335, p => False), (a => 175, b => 239, p => False), (a => 159, b => 223, p => False), (a => 287, b => 351, p => False), (a => 288, b => 320, p => False), (a => 0  , b => 319, p => True ), (a => 1  , b => 318, p => True ), (a => 62 , b => 317, p => True ), (a => 63 , b => 316, p => True ), (a => 64 , b => 315, p => True ), (a => 65 , b => 314, p => True ), (a => 66 , b => 313, p => True ), (a => 67 , b => 312, p => True ), (a => 68 , b => 311, p => True ), (a => 69 , b => 310, p => True ), (a => 70 , b => 309, p => True ), (a => 71 , b => 308, p => True ), (a => 72 , b => 307, p => True ), (a => 73 , b => 306, p => True ), (a => 74 , b => 305, p => True ), (a => 75 , b => 304, p => True ), (a => 76 , b => 303, p => True ), (a => 77 , b => 302, p => True ), (a => 78 , b => 301, p => True ), (a => 79 , b => 300, p => True ), (a => 80 , b => 299, p => True ), (a => 81 , b => 298, p => True ), (a => 82 , b => 297, p => True ), (a => 83 , b => 296, p => True ), (a => 84 , b => 295, p => True ), (a => 85 , b => 294, p => True ), (a => 86 , b => 293, p => True ), (a => 87 , b => 292, p => True ), (a => 88 , b => 291, p => True ), (a => 89 , b => 290, p => True ), (a => 90 , b => 289, p => True ), (a => 91 , b => 256, p => True ), (a => 92 , b => 255, p => True ), (a => 93 , b => 192, p => True ), (a => 94 , b => 191, p => True ), (a => 95 , b => 128, p => True ), (a => 96 , b => 127, p => True ), (a => 97 , b => 126, p => True ), (a => 98 , b => 125, p => True ), (a => 99 , b => 124, p => True ), (a => 100, b => 123, p => True ), (a => 101, b => 122, p => True ), (a => 102, b => 121, p => True ), (a => 103, b => 120, p => True ), (a => 104, b => 119, p => True ), (a => 105, b => 118, p => True ), (a => 106, b => 117, p => True ), (a => 107, b => 116, p => True ), (a => 108, b => 115, p => True ), (a => 109, b => 114, p => True ), (a => 110, b => 113, p => True ), (a => 111, b => 112, p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 31 , b => 32 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 47 , b => 48 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 160, b => 192, p => False), (a => 176, b => 208, p => False), (a => 304, b => 336, p => False), (a => 168, b => 200, p => False), (a => 296, b => 328, p => False), (a => 184, b => 216, p => False), (a => 312, b => 344, p => False), (a => 164, b => 196, p => False), (a => 292, b => 324, p => False), (a => 180, b => 212, p => False), (a => 308, b => 340, p => False), (a => 172, b => 204, p => False), (a => 300, b => 332, p => False), (a => 188, b => 220, p => False), (a => 316, b => 348, p => False), (a => 162, b => 194, p => False), (a => 290, b => 322, p => False), (a => 178, b => 210, p => False), (a => 306, b => 338, p => False), (a => 170, b => 202, p => False), (a => 298, b => 330, p => False), (a => 186, b => 218, p => False), (a => 314, b => 346, p => False), (a => 166, b => 198, p => False), (a => 294, b => 326, p => False), (a => 182, b => 214, p => False), (a => 310, b => 342, p => False), (a => 174, b => 206, p => False), (a => 302, b => 334, p => False), (a => 190, b => 222, p => False), (a => 318, b => 350, p => False), (a => 161, b => 193, p => False), (a => 289, b => 321, p => False), (a => 177, b => 209, p => False), (a => 305, b => 337, p => False), (a => 169, b => 201, p => False), (a => 297, b => 329, p => False), (a => 185, b => 217, p => False), (a => 313, b => 345, p => False), (a => 165, b => 197, p => False), (a => 293, b => 325, p => False), (a => 181, b => 213, p => False), (a => 309, b => 341, p => False), (a => 173, b => 205, p => False), (a => 301, b => 333, p => False), (a => 189, b => 221, p => False), (a => 317, b => 349, p => False), (a => 163, b => 195, p => False), (a => 291, b => 323, p => False), (a => 179, b => 211, p => False), (a => 307, b => 339, p => False), (a => 171, b => 203, p => False), (a => 299, b => 331, p => False), (a => 187, b => 219, p => False), (a => 315, b => 347, p => False), (a => 167, b => 199, p => False), (a => 295, b => 327, p => False), (a => 183, b => 215, p => False), (a => 311, b => 343, p => False), (a => 175, b => 207, p => False), (a => 303, b => 335, p => False), (a => 191, b => 223, p => False), (a => 319, b => 351, p => False), (a => 272, b => 288, p => False), (a => 0  , b => 320, p => True ), (a => 63 , b => 287, p => True ), (a => 64 , b => 286, p => True ), (a => 65 , b => 285, p => True ), (a => 66 , b => 284, p => True ), (a => 67 , b => 283, p => True ), (a => 68 , b => 282, p => True ), (a => 69 , b => 281, p => True ), (a => 70 , b => 280, p => True ), (a => 71 , b => 279, p => True ), (a => 72 , b => 278, p => True ), (a => 73 , b => 277, p => True ), (a => 74 , b => 276, p => True ), (a => 75 , b => 275, p => True ), (a => 76 , b => 274, p => True ), (a => 77 , b => 273, p => True ), (a => 78 , b => 271, p => True ), (a => 79 , b => 270, p => True ), (a => 80 , b => 269, p => True ), (a => 81 , b => 268, p => True ), (a => 82 , b => 267, p => True ), (a => 83 , b => 266, p => True ), (a => 84 , b => 265, p => True ), (a => 85 , b => 264, p => True ), (a => 86 , b => 263, p => True ), (a => 87 , b => 262, p => True ), (a => 88 , b => 261, p => True ), (a => 89 , b => 260, p => True ), (a => 90 , b => 259, p => True ), (a => 91 , b => 258, p => True ), (a => 92 , b => 257, p => True ), (a => 93 , b => 256, p => True ), (a => 94 , b => 255, p => True ), (a => 95 , b => 254, p => True ), (a => 96 , b => 253, p => True ), (a => 97 , b => 252, p => True ), (a => 98 , b => 251, p => True ), (a => 99 , b => 250, p => True ), (a => 100, b => 249, p => True ), (a => 101, b => 248, p => True ), (a => 102, b => 247, p => True ), (a => 103, b => 246, p => True ), (a => 104, b => 245, p => True ), (a => 105, b => 244, p => True ), (a => 106, b => 243, p => True ), (a => 107, b => 242, p => True ), (a => 108, b => 241, p => True ), (a => 109, b => 240, p => True ), (a => 110, b => 239, p => True ), (a => 111, b => 238, p => True ), (a => 112, b => 237, p => True ), (a => 113, b => 236, p => True ), (a => 114, b => 235, p => True ), (a => 115, b => 234, p => True ), (a => 116, b => 233, p => True ), (a => 117, b => 232, p => True ), (a => 118, b => 231, p => True ), (a => 119, b => 230, p => True ), (a => 120, b => 229, p => True ), (a => 121, b => 228, p => True ), (a => 122, b => 227, p => True ), (a => 123, b => 226, p => True ), (a => 124, b => 225, p => True ), (a => 125, b => 224, p => True ), (a => 126, b => 159, p => True ), (a => 127, b => 158, p => True ), (a => 128, b => 157, p => True ), (a => 129, b => 156, p => True ), (a => 130, b => 155, p => True ), (a => 131, b => 154, p => True ), (a => 132, b => 153, p => True ), (a => 133, b => 152, p => True ), (a => 134, b => 151, p => True ), (a => 135, b => 150, p => True ), (a => 136, b => 149, p => True ), (a => 137, b => 148, p => True ), (a => 138, b => 147, p => True ), (a => 139, b => 146, p => True ), (a => 140, b => 145, p => True ), (a => 141, b => 144, p => True ), (a => 142, b => 143, p => True )),
                    ((a => 32 , b => 96 , p => False), (a => 16 , b => 80 , p => False), (a => 48 , b => 112, p => False), (a => 8  , b => 72 , p => False), (a => 40 , b => 104, p => False), (a => 24 , b => 88 , p => False), (a => 56 , b => 120, p => False), (a => 4  , b => 68 , p => False), (a => 36 , b => 100, p => False), (a => 20 , b => 84 , p => False), (a => 52 , b => 116, p => False), (a => 12 , b => 76 , p => False), (a => 44 , b => 108, p => False), (a => 28 , b => 92 , p => False), (a => 60 , b => 124, p => False), (a => 2  , b => 66 , p => False), (a => 34 , b => 98 , p => False), (a => 18 , b => 82 , p => False), (a => 50 , b => 114, p => False), (a => 10 , b => 74 , p => False), (a => 42 , b => 106, p => False), (a => 26 , b => 90 , p => False), (a => 58 , b => 122, p => False), (a => 6  , b => 70 , p => False), (a => 38 , b => 102, p => False), (a => 22 , b => 86 , p => False), (a => 54 , b => 118, p => False), (a => 14 , b => 78 , p => False), (a => 46 , b => 110, p => False), (a => 30 , b => 94 , p => False), (a => 62 , b => 126, p => False), (a => 1  , b => 65 , p => False), (a => 33 , b => 97 , p => False), (a => 17 , b => 81 , p => False), (a => 49 , b => 113, p => False), (a => 9  , b => 73 , p => False), (a => 41 , b => 105, p => False), (a => 25 , b => 89 , p => False), (a => 57 , b => 121, p => False), (a => 5  , b => 69 , p => False), (a => 37 , b => 101, p => False), (a => 21 , b => 85 , p => False), (a => 53 , b => 117, p => False), (a => 13 , b => 77 , p => False), (a => 45 , b => 109, p => False), (a => 29 , b => 93 , p => False), (a => 61 , b => 125, p => False), (a => 3  , b => 67 , p => False), (a => 35 , b => 99 , p => False), (a => 19 , b => 83 , p => False), (a => 51 , b => 115, p => False), (a => 11 , b => 75 , p => False), (a => 43 , b => 107, p => False), (a => 27 , b => 91 , p => False), (a => 59 , b => 123, p => False), (a => 7  , b => 71 , p => False), (a => 39 , b => 103, p => False), (a => 23 , b => 87 , p => False), (a => 55 , b => 119, p => False), (a => 15 , b => 79 , p => False), (a => 47 , b => 111, p => False), (a => 31 , b => 95 , p => False), (a => 144, b => 160, p => False), (a => 176, b => 192, p => False), (a => 208, b => 224, p => False), (a => 304, b => 320, p => False), (a => 152, b => 168, p => False), (a => 184, b => 200, p => False), (a => 216, b => 232, p => False), (a => 280, b => 296, p => False), (a => 312, b => 328, p => False), (a => 148, b => 164, p => False), (a => 180, b => 196, p => False), (a => 212, b => 228, p => False), (a => 276, b => 292, p => False), (a => 308, b => 324, p => False), (a => 156, b => 172, p => False), (a => 188, b => 204, p => False), (a => 220, b => 236, p => False), (a => 284, b => 300, p => False), (a => 316, b => 332, p => False), (a => 146, b => 162, p => False), (a => 178, b => 194, p => False), (a => 210, b => 226, p => False), (a => 274, b => 290, p => False), (a => 306, b => 322, p => False), (a => 154, b => 170, p => False), (a => 186, b => 202, p => False), (a => 218, b => 234, p => False), (a => 282, b => 298, p => False), (a => 314, b => 330, p => False), (a => 150, b => 166, p => False), (a => 182, b => 198, p => False), (a => 214, b => 230, p => False), (a => 278, b => 294, p => False), (a => 310, b => 326, p => False), (a => 158, b => 174, p => False), (a => 190, b => 206, p => False), (a => 222, b => 238, p => False), (a => 286, b => 302, p => False), (a => 318, b => 334, p => False), (a => 145, b => 161, p => False), (a => 177, b => 193, p => False), (a => 209, b => 225, p => False), (a => 273, b => 289, p => False), (a => 305, b => 321, p => False), (a => 153, b => 169, p => False), (a => 185, b => 201, p => False), (a => 217, b => 233, p => False), (a => 281, b => 297, p => False), (a => 313, b => 329, p => False), (a => 149, b => 165, p => False), (a => 181, b => 197, p => False), (a => 213, b => 229, p => False), (a => 277, b => 293, p => False), (a => 309, b => 325, p => False), (a => 157, b => 173, p => False), (a => 189, b => 205, p => False), (a => 221, b => 237, p => False), (a => 285, b => 301, p => False), (a => 317, b => 333, p => False), (a => 147, b => 163, p => False), (a => 179, b => 195, p => False), (a => 211, b => 227, p => False), (a => 275, b => 291, p => False), (a => 307, b => 323, p => False), (a => 155, b => 171, p => False), (a => 187, b => 203, p => False), (a => 219, b => 235, p => False), (a => 283, b => 299, p => False), (a => 315, b => 331, p => False), (a => 151, b => 167, p => False), (a => 183, b => 199, p => False), (a => 215, b => 231, p => False), (a => 279, b => 295, p => False), (a => 311, b => 327, p => False), (a => 159, b => 175, p => False), (a => 191, b => 207, p => False), (a => 223, b => 239, p => False), (a => 287, b => 303, p => False), (a => 319, b => 335, p => False), (a => 264, b => 272, p => False), (a => 0  , b => 351, p => True ), (a => 63 , b => 350, p => True ), (a => 64 , b => 349, p => True ), (a => 127, b => 348, p => True ), (a => 128, b => 347, p => True ), (a => 129, b => 346, p => True ), (a => 130, b => 345, p => True ), (a => 131, b => 344, p => True ), (a => 132, b => 343, p => True ), (a => 133, b => 342, p => True ), (a => 134, b => 341, p => True ), (a => 135, b => 340, p => True ), (a => 136, b => 339, p => True ), (a => 137, b => 338, p => True ), (a => 138, b => 337, p => True ), (a => 139, b => 336, p => True ), (a => 140, b => 288, p => True ), (a => 141, b => 271, p => True ), (a => 142, b => 270, p => True ), (a => 143, b => 269, p => True ), (a => 240, b => 268, p => True ), (a => 241, b => 267, p => True ), (a => 242, b => 266, p => True ), (a => 243, b => 265, p => True ), (a => 244, b => 263, p => True ), (a => 245, b => 262, p => True ), (a => 246, b => 261, p => True ), (a => 247, b => 260, p => True ), (a => 248, b => 259, p => True ), (a => 249, b => 258, p => True ), (a => 250, b => 257, p => True ), (a => 251, b => 256, p => True ), (a => 252, b => 255, p => True ), (a => 253, b => 254, p => True )),
                    ((a => 32 , b => 64 , p => False), (a => 48 , b => 80 , p => False), (a => 40 , b => 72 , p => False), (a => 56 , b => 88 , p => False), (a => 36 , b => 68 , p => False), (a => 52 , b => 84 , p => False), (a => 44 , b => 76 , p => False), (a => 60 , b => 92 , p => False), (a => 34 , b => 66 , p => False), (a => 50 , b => 82 , p => False), (a => 42 , b => 74 , p => False), (a => 58 , b => 90 , p => False), (a => 38 , b => 70 , p => False), (a => 54 , b => 86 , p => False), (a => 46 , b => 78 , p => False), (a => 62 , b => 94 , p => False), (a => 33 , b => 65 , p => False), (a => 49 , b => 81 , p => False), (a => 41 , b => 73 , p => False), (a => 57 , b => 89 , p => False), (a => 37 , b => 69 , p => False), (a => 53 , b => 85 , p => False), (a => 45 , b => 77 , p => False), (a => 61 , b => 93 , p => False), (a => 35 , b => 67 , p => False), (a => 51 , b => 83 , p => False), (a => 43 , b => 75 , p => False), (a => 59 , b => 91 , p => False), (a => 39 , b => 71 , p => False), (a => 55 , b => 87 , p => False), (a => 47 , b => 79 , p => False), (a => 63 , b => 95 , p => False), (a => 136, b => 144, p => False), (a => 152, b => 160, p => False), (a => 168, b => 176, p => False), (a => 184, b => 192, p => False), (a => 200, b => 208, p => False), (a => 216, b => 224, p => False), (a => 232, b => 240, p => False), (a => 280, b => 288, p => False), (a => 296, b => 304, p => False), (a => 312, b => 320, p => False), (a => 328, b => 336, p => False), (a => 140, b => 148, p => False), (a => 156, b => 164, p => False), (a => 172, b => 180, p => False), (a => 188, b => 196, p => False), (a => 204, b => 212, p => False), (a => 220, b => 228, p => False), (a => 236, b => 244, p => False), (a => 268, b => 276, p => False), (a => 284, b => 292, p => False), (a => 300, b => 308, p => False), (a => 316, b => 324, p => False), (a => 332, b => 340, p => False), (a => 138, b => 146, p => False), (a => 154, b => 162, p => False), (a => 170, b => 178, p => False), (a => 186, b => 194, p => False), (a => 202, b => 210, p => False), (a => 218, b => 226, p => False), (a => 234, b => 242, p => False), (a => 266, b => 274, p => False), (a => 282, b => 290, p => False), (a => 298, b => 306, p => False), (a => 314, b => 322, p => False), (a => 330, b => 338, p => False), (a => 142, b => 150, p => False), (a => 158, b => 166, p => False), (a => 174, b => 182, p => False), (a => 190, b => 198, p => False), (a => 206, b => 214, p => False), (a => 222, b => 230, p => False), (a => 238, b => 246, p => False), (a => 270, b => 278, p => False), (a => 286, b => 294, p => False), (a => 302, b => 310, p => False), (a => 318, b => 326, p => False), (a => 334, b => 342, p => False), (a => 137, b => 145, p => False), (a => 153, b => 161, p => False), (a => 169, b => 177, p => False), (a => 185, b => 193, p => False), (a => 201, b => 209, p => False), (a => 217, b => 225, p => False), (a => 233, b => 241, p => False), (a => 265, b => 273, p => False), (a => 281, b => 289, p => False), (a => 297, b => 305, p => False), (a => 313, b => 321, p => False), (a => 329, b => 337, p => False), (a => 141, b => 149, p => False), (a => 157, b => 165, p => False), (a => 173, b => 181, p => False), (a => 189, b => 197, p => False), (a => 205, b => 213, p => False), (a => 221, b => 229, p => False), (a => 237, b => 245, p => False), (a => 269, b => 277, p => False), (a => 285, b => 293, p => False), (a => 301, b => 309, p => False), (a => 317, b => 325, p => False), (a => 333, b => 341, p => False), (a => 139, b => 147, p => False), (a => 155, b => 163, p => False), (a => 171, b => 179, p => False), (a => 187, b => 195, p => False), (a => 203, b => 211, p => False), (a => 219, b => 227, p => False), (a => 235, b => 243, p => False), (a => 267, b => 275, p => False), (a => 283, b => 291, p => False), (a => 299, b => 307, p => False), (a => 315, b => 323, p => False), (a => 331, b => 339, p => False), (a => 143, b => 151, p => False), (a => 159, b => 167, p => False), (a => 175, b => 183, p => False), (a => 191, b => 199, p => False), (a => 207, b => 215, p => False), (a => 223, b => 231, p => False), (a => 239, b => 247, p => False), (a => 271, b => 279, p => False), (a => 287, b => 295, p => False), (a => 303, b => 311, p => False), (a => 319, b => 327, p => False), (a => 335, b => 343, p => False), (a => 260, b => 264, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 272, p => True ), (a => 9  , b => 263, p => True ), (a => 10 , b => 262, p => True ), (a => 11 , b => 261, p => True ), (a => 12 , b => 259, p => True ), (a => 13 , b => 258, p => True ), (a => 14 , b => 257, p => True ), (a => 15 , b => 256, p => True ), (a => 16 , b => 255, p => True ), (a => 17 , b => 254, p => True ), (a => 18 , b => 253, p => True ), (a => 19 , b => 252, p => True ), (a => 20 , b => 251, p => True ), (a => 21 , b => 250, p => True ), (a => 22 , b => 249, p => True ), (a => 23 , b => 248, p => True ), (a => 24 , b => 135, p => True ), (a => 25 , b => 134, p => True ), (a => 26 , b => 133, p => True ), (a => 27 , b => 132, p => True ), (a => 28 , b => 131, p => True ), (a => 29 , b => 130, p => True ), (a => 30 , b => 129, p => True ), (a => 31 , b => 128, p => True ), (a => 96 , b => 127, p => True ), (a => 97 , b => 126, p => True ), (a => 98 , b => 125, p => True ), (a => 99 , b => 124, p => True ), (a => 100, b => 123, p => True ), (a => 101, b => 122, p => True ), (a => 102, b => 121, p => True ), (a => 103, b => 120, p => True ), (a => 104, b => 119, p => True ), (a => 105, b => 118, p => True ), (a => 106, b => 117, p => True ), (a => 107, b => 116, p => True ), (a => 108, b => 115, p => True ), (a => 109, b => 114, p => True ), (a => 110, b => 113, p => True ), (a => 111, b => 112, p => True )),
                    ((a => 16 , b => 32 , p => False), (a => 48 , b => 64 , p => False), (a => 80 , b => 96 , p => False), (a => 24 , b => 40 , p => False), (a => 56 , b => 72 , p => False), (a => 88 , b => 104, p => False), (a => 20 , b => 36 , p => False), (a => 52 , b => 68 , p => False), (a => 84 , b => 100, p => False), (a => 28 , b => 44 , p => False), (a => 60 , b => 76 , p => False), (a => 92 , b => 108, p => False), (a => 18 , b => 34 , p => False), (a => 50 , b => 66 , p => False), (a => 82 , b => 98 , p => False), (a => 26 , b => 42 , p => False), (a => 58 , b => 74 , p => False), (a => 90 , b => 106, p => False), (a => 22 , b => 38 , p => False), (a => 54 , b => 70 , p => False), (a => 86 , b => 102, p => False), (a => 30 , b => 46 , p => False), (a => 62 , b => 78 , p => False), (a => 94 , b => 110, p => False), (a => 17 , b => 33 , p => False), (a => 49 , b => 65 , p => False), (a => 81 , b => 97 , p => False), (a => 25 , b => 41 , p => False), (a => 57 , b => 73 , p => False), (a => 89 , b => 105, p => False), (a => 21 , b => 37 , p => False), (a => 53 , b => 69 , p => False), (a => 85 , b => 101, p => False), (a => 29 , b => 45 , p => False), (a => 61 , b => 77 , p => False), (a => 93 , b => 109, p => False), (a => 19 , b => 35 , p => False), (a => 51 , b => 67 , p => False), (a => 83 , b => 99 , p => False), (a => 27 , b => 43 , p => False), (a => 59 , b => 75 , p => False), (a => 91 , b => 107, p => False), (a => 23 , b => 39 , p => False), (a => 55 , b => 71 , p => False), (a => 87 , b => 103, p => False), (a => 31 , b => 47 , p => False), (a => 63 , b => 79 , p => False), (a => 95 , b => 111, p => False), (a => 132, b => 136, p => False), (a => 140, b => 144, p => False), (a => 148, b => 152, p => False), (a => 156, b => 160, p => False), (a => 164, b => 168, p => False), (a => 172, b => 176, p => False), (a => 180, b => 184, p => False), (a => 188, b => 192, p => False), (a => 196, b => 200, p => False), (a => 204, b => 208, p => False), (a => 212, b => 216, p => False), (a => 220, b => 224, p => False), (a => 228, b => 232, p => False), (a => 236, b => 240, p => False), (a => 244, b => 248, p => False), (a => 268, b => 272, p => False), (a => 276, b => 280, p => False), (a => 284, b => 288, p => False), (a => 292, b => 296, p => False), (a => 300, b => 304, p => False), (a => 308, b => 312, p => False), (a => 316, b => 320, p => False), (a => 324, b => 328, p => False), (a => 332, b => 336, p => False), (a => 340, b => 344, p => False), (a => 134, b => 138, p => False), (a => 142, b => 146, p => False), (a => 150, b => 154, p => False), (a => 158, b => 162, p => False), (a => 166, b => 170, p => False), (a => 174, b => 178, p => False), (a => 182, b => 186, p => False), (a => 190, b => 194, p => False), (a => 198, b => 202, p => False), (a => 206, b => 210, p => False), (a => 214, b => 218, p => False), (a => 222, b => 226, p => False), (a => 230, b => 234, p => False), (a => 238, b => 242, p => False), (a => 246, b => 250, p => False), (a => 262, b => 266, p => False), (a => 270, b => 274, p => False), (a => 278, b => 282, p => False), (a => 286, b => 290, p => False), (a => 294, b => 298, p => False), (a => 302, b => 306, p => False), (a => 310, b => 314, p => False), (a => 318, b => 322, p => False), (a => 326, b => 330, p => False), (a => 334, b => 338, p => False), (a => 342, b => 346, p => False), (a => 133, b => 137, p => False), (a => 141, b => 145, p => False), (a => 149, b => 153, p => False), (a => 157, b => 161, p => False), (a => 165, b => 169, p => False), (a => 173, b => 177, p => False), (a => 181, b => 185, p => False), (a => 189, b => 193, p => False), (a => 197, b => 201, p => False), (a => 205, b => 209, p => False), (a => 213, b => 217, p => False), (a => 221, b => 225, p => False), (a => 229, b => 233, p => False), (a => 237, b => 241, p => False), (a => 245, b => 249, p => False), (a => 261, b => 265, p => False), (a => 269, b => 273, p => False), (a => 277, b => 281, p => False), (a => 285, b => 289, p => False), (a => 293, b => 297, p => False), (a => 301, b => 305, p => False), (a => 309, b => 313, p => False), (a => 317, b => 321, p => False), (a => 325, b => 329, p => False), (a => 333, b => 337, p => False), (a => 341, b => 345, p => False), (a => 135, b => 139, p => False), (a => 143, b => 147, p => False), (a => 151, b => 155, p => False), (a => 159, b => 163, p => False), (a => 167, b => 171, p => False), (a => 175, b => 179, p => False), (a => 183, b => 187, p => False), (a => 191, b => 195, p => False), (a => 199, b => 203, p => False), (a => 207, b => 211, p => False), (a => 215, b => 219, p => False), (a => 223, b => 227, p => False), (a => 231, b => 235, p => False), (a => 239, b => 243, p => False), (a => 247, b => 251, p => False), (a => 263, b => 267, p => False), (a => 271, b => 275, p => False), (a => 279, b => 283, p => False), (a => 287, b => 291, p => False), (a => 295, b => 299, p => False), (a => 303, b => 307, p => False), (a => 311, b => 315, p => False), (a => 319, b => 323, p => False), (a => 327, b => 331, p => False), (a => 335, b => 339, p => False), (a => 343, b => 347, p => False), (a => 258, b => 260, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 264, p => True ), (a => 5  , b => 259, p => True ), (a => 6  , b => 257, p => True ), (a => 7  , b => 256, p => True ), (a => 8  , b => 255, p => True ), (a => 9  , b => 254, p => True ), (a => 10 , b => 253, p => True ), (a => 11 , b => 252, p => True ), (a => 12 , b => 131, p => True ), (a => 13 , b => 130, p => True ), (a => 14 , b => 129, p => True ), (a => 15 , b => 128, p => True ), (a => 112, b => 127, p => True ), (a => 113, b => 126, p => True ), (a => 114, b => 125, p => True ), (a => 115, b => 124, p => True ), (a => 116, b => 123, p => True ), (a => 117, b => 122, p => True ), (a => 118, b => 121, p => True ), (a => 119, b => 120, p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 24 , b => 32 , p => False), (a => 40 , b => 48 , p => False), (a => 56 , b => 64 , p => False), (a => 72 , b => 80 , p => False), (a => 88 , b => 96 , p => False), (a => 104, b => 112, p => False), (a => 12 , b => 20 , p => False), (a => 28 , b => 36 , p => False), (a => 44 , b => 52 , p => False), (a => 60 , b => 68 , p => False), (a => 76 , b => 84 , p => False), (a => 92 , b => 100, p => False), (a => 108, b => 116, p => False), (a => 10 , b => 18 , p => False), (a => 26 , b => 34 , p => False), (a => 42 , b => 50 , p => False), (a => 58 , b => 66 , p => False), (a => 74 , b => 82 , p => False), (a => 90 , b => 98 , p => False), (a => 106, b => 114, p => False), (a => 14 , b => 22 , p => False), (a => 30 , b => 38 , p => False), (a => 46 , b => 54 , p => False), (a => 62 , b => 70 , p => False), (a => 78 , b => 86 , p => False), (a => 94 , b => 102, p => False), (a => 110, b => 118, p => False), (a => 9  , b => 17 , p => False), (a => 25 , b => 33 , p => False), (a => 41 , b => 49 , p => False), (a => 57 , b => 65 , p => False), (a => 73 , b => 81 , p => False), (a => 89 , b => 97 , p => False), (a => 105, b => 113, p => False), (a => 13 , b => 21 , p => False), (a => 29 , b => 37 , p => False), (a => 45 , b => 53 , p => False), (a => 61 , b => 69 , p => False), (a => 77 , b => 85 , p => False), (a => 93 , b => 101, p => False), (a => 109, b => 117, p => False), (a => 11 , b => 19 , p => False), (a => 27 , b => 35 , p => False), (a => 43 , b => 51 , p => False), (a => 59 , b => 67 , p => False), (a => 75 , b => 83 , p => False), (a => 91 , b => 99 , p => False), (a => 107, b => 115, p => False), (a => 15 , b => 23 , p => False), (a => 31 , b => 39 , p => False), (a => 47 , b => 55 , p => False), (a => 63 , b => 71 , p => False), (a => 79 , b => 87 , p => False), (a => 95 , b => 103, p => False), (a => 111, b => 119, p => False), (a => 130, b => 132, p => False), (a => 134, b => 136, p => False), (a => 138, b => 140, p => False), (a => 142, b => 144, p => False), (a => 146, b => 148, p => False), (a => 150, b => 152, p => False), (a => 154, b => 156, p => False), (a => 158, b => 160, p => False), (a => 162, b => 164, p => False), (a => 166, b => 168, p => False), (a => 170, b => 172, p => False), (a => 174, b => 176, p => False), (a => 178, b => 180, p => False), (a => 182, b => 184, p => False), (a => 186, b => 188, p => False), (a => 190, b => 192, p => False), (a => 194, b => 196, p => False), (a => 198, b => 200, p => False), (a => 202, b => 204, p => False), (a => 206, b => 208, p => False), (a => 210, b => 212, p => False), (a => 214, b => 216, p => False), (a => 218, b => 220, p => False), (a => 222, b => 224, p => False), (a => 226, b => 228, p => False), (a => 230, b => 232, p => False), (a => 234, b => 236, p => False), (a => 238, b => 240, p => False), (a => 242, b => 244, p => False), (a => 246, b => 248, p => False), (a => 250, b => 252, p => False), (a => 262, b => 264, p => False), (a => 266, b => 268, p => False), (a => 270, b => 272, p => False), (a => 274, b => 276, p => False), (a => 278, b => 280, p => False), (a => 282, b => 284, p => False), (a => 286, b => 288, p => False), (a => 290, b => 292, p => False), (a => 294, b => 296, p => False), (a => 298, b => 300, p => False), (a => 302, b => 304, p => False), (a => 306, b => 308, p => False), (a => 310, b => 312, p => False), (a => 314, b => 316, p => False), (a => 318, b => 320, p => False), (a => 322, b => 324, p => False), (a => 326, b => 328, p => False), (a => 330, b => 332, p => False), (a => 334, b => 336, p => False), (a => 338, b => 340, p => False), (a => 342, b => 344, p => False), (a => 346, b => 348, p => False), (a => 131, b => 133, p => False), (a => 135, b => 137, p => False), (a => 139, b => 141, p => False), (a => 143, b => 145, p => False), (a => 147, b => 149, p => False), (a => 151, b => 153, p => False), (a => 155, b => 157, p => False), (a => 159, b => 161, p => False), (a => 163, b => 165, p => False), (a => 167, b => 169, p => False), (a => 171, b => 173, p => False), (a => 175, b => 177, p => False), (a => 179, b => 181, p => False), (a => 183, b => 185, p => False), (a => 187, b => 189, p => False), (a => 191, b => 193, p => False), (a => 195, b => 197, p => False), (a => 199, b => 201, p => False), (a => 203, b => 205, p => False), (a => 207, b => 209, p => False), (a => 211, b => 213, p => False), (a => 215, b => 217, p => False), (a => 219, b => 221, p => False), (a => 223, b => 225, p => False), (a => 227, b => 229, p => False), (a => 231, b => 233, p => False), (a => 235, b => 237, p => False), (a => 239, b => 241, p => False), (a => 243, b => 245, p => False), (a => 247, b => 249, p => False), (a => 251, b => 253, p => False), (a => 259, b => 261, p => False), (a => 263, b => 265, p => False), (a => 267, b => 269, p => False), (a => 271, b => 273, p => False), (a => 275, b => 277, p => False), (a => 279, b => 281, p => False), (a => 283, b => 285, p => False), (a => 287, b => 289, p => False), (a => 291, b => 293, p => False), (a => 295, b => 297, p => False), (a => 299, b => 301, p => False), (a => 303, b => 305, p => False), (a => 307, b => 309, p => False), (a => 311, b => 313, p => False), (a => 315, b => 317, p => False), (a => 319, b => 321, p => False), (a => 323, b => 325, p => False), (a => 327, b => 329, p => False), (a => 331, b => 333, p => False), (a => 335, b => 337, p => False), (a => 339, b => 341, p => False), (a => 343, b => 345, p => False), (a => 347, b => 349, p => False), (a => 257, b => 258, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 260, p => True ), (a => 3  , b => 256, p => True ), (a => 4  , b => 255, p => True ), (a => 5  , b => 254, p => True ), (a => 6  , b => 129, p => True ), (a => 7  , b => 128, p => True ), (a => 120, b => 127, p => True ), (a => 121, b => 126, p => True ), (a => 122, b => 125, p => True ), (a => 123, b => 124, p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 28 , b => 32 , p => False), (a => 36 , b => 40 , p => False), (a => 44 , b => 48 , p => False), (a => 52 , b => 56 , p => False), (a => 60 , b => 64 , p => False), (a => 68 , b => 72 , p => False), (a => 76 , b => 80 , p => False), (a => 84 , b => 88 , p => False), (a => 92 , b => 96 , p => False), (a => 100, b => 104, p => False), (a => 108, b => 112, p => False), (a => 116, b => 120, p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 30 , b => 34 , p => False), (a => 38 , b => 42 , p => False), (a => 46 , b => 50 , p => False), (a => 54 , b => 58 , p => False), (a => 62 , b => 66 , p => False), (a => 70 , b => 74 , p => False), (a => 78 , b => 82 , p => False), (a => 86 , b => 90 , p => False), (a => 94 , b => 98 , p => False), (a => 102, b => 106, p => False), (a => 110, b => 114, p => False), (a => 118, b => 122, p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 29 , b => 33 , p => False), (a => 37 , b => 41 , p => False), (a => 45 , b => 49 , p => False), (a => 53 , b => 57 , p => False), (a => 61 , b => 65 , p => False), (a => 69 , b => 73 , p => False), (a => 77 , b => 81 , p => False), (a => 85 , b => 89 , p => False), (a => 93 , b => 97 , p => False), (a => 101, b => 105, p => False), (a => 109, b => 113, p => False), (a => 117, b => 121, p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 31 , b => 35 , p => False), (a => 39 , b => 43 , p => False), (a => 47 , b => 51 , p => False), (a => 55 , b => 59 , p => False), (a => 63 , b => 67 , p => False), (a => 71 , b => 75 , p => False), (a => 79 , b => 83 , p => False), (a => 87 , b => 91 , p => False), (a => 95 , b => 99 , p => False), (a => 103, b => 107, p => False), (a => 111, b => 115, p => False), (a => 119, b => 123, p => False), (a => 129, b => 130, p => False), (a => 131, b => 132, p => False), (a => 133, b => 134, p => False), (a => 135, b => 136, p => False), (a => 137, b => 138, p => False), (a => 139, b => 140, p => False), (a => 141, b => 142, p => False), (a => 143, b => 144, p => False), (a => 145, b => 146, p => False), (a => 147, b => 148, p => False), (a => 149, b => 150, p => False), (a => 151, b => 152, p => False), (a => 153, b => 154, p => False), (a => 155, b => 156, p => False), (a => 157, b => 158, p => False), (a => 159, b => 160, p => False), (a => 161, b => 162, p => False), (a => 163, b => 164, p => False), (a => 165, b => 166, p => False), (a => 167, b => 168, p => False), (a => 169, b => 170, p => False), (a => 171, b => 172, p => False), (a => 173, b => 174, p => False), (a => 175, b => 176, p => False), (a => 177, b => 178, p => False), (a => 179, b => 180, p => False), (a => 181, b => 182, p => False), (a => 183, b => 184, p => False), (a => 185, b => 186, p => False), (a => 187, b => 188, p => False), (a => 189, b => 190, p => False), (a => 191, b => 192, p => False), (a => 193, b => 194, p => False), (a => 195, b => 196, p => False), (a => 197, b => 198, p => False), (a => 199, b => 200, p => False), (a => 201, b => 202, p => False), (a => 203, b => 204, p => False), (a => 205, b => 206, p => False), (a => 207, b => 208, p => False), (a => 209, b => 210, p => False), (a => 211, b => 212, p => False), (a => 213, b => 214, p => False), (a => 215, b => 216, p => False), (a => 217, b => 218, p => False), (a => 219, b => 220, p => False), (a => 221, b => 222, p => False), (a => 223, b => 224, p => False), (a => 225, b => 226, p => False), (a => 227, b => 228, p => False), (a => 229, b => 230, p => False), (a => 231, b => 232, p => False), (a => 233, b => 234, p => False), (a => 235, b => 236, p => False), (a => 237, b => 238, p => False), (a => 239, b => 240, p => False), (a => 241, b => 242, p => False), (a => 243, b => 244, p => False), (a => 245, b => 246, p => False), (a => 247, b => 248, p => False), (a => 249, b => 250, p => False), (a => 251, b => 252, p => False), (a => 253, b => 254, p => False), (a => 259, b => 260, p => False), (a => 261, b => 262, p => False), (a => 263, b => 264, p => False), (a => 265, b => 266, p => False), (a => 267, b => 268, p => False), (a => 269, b => 270, p => False), (a => 271, b => 272, p => False), (a => 273, b => 274, p => False), (a => 275, b => 276, p => False), (a => 277, b => 278, p => False), (a => 279, b => 280, p => False), (a => 281, b => 282, p => False), (a => 283, b => 284, p => False), (a => 285, b => 286, p => False), (a => 287, b => 288, p => False), (a => 289, b => 290, p => False), (a => 291, b => 292, p => False), (a => 293, b => 294, p => False), (a => 295, b => 296, p => False), (a => 297, b => 298, p => False), (a => 299, b => 300, p => False), (a => 301, b => 302, p => False), (a => 303, b => 304, p => False), (a => 305, b => 306, p => False), (a => 307, b => 308, p => False), (a => 309, b => 310, p => False), (a => 311, b => 312, p => False), (a => 313, b => 314, p => False), (a => 315, b => 316, p => False), (a => 317, b => 318, p => False), (a => 319, b => 320, p => False), (a => 321, b => 322, p => False), (a => 323, b => 324, p => False), (a => 325, b => 326, p => False), (a => 327, b => 328, p => False), (a => 329, b => 330, p => False), (a => 331, b => 332, p => False), (a => 333, b => 334, p => False), (a => 335, b => 336, p => False), (a => 337, b => 338, p => False), (a => 339, b => 340, p => False), (a => 341, b => 342, p => False), (a => 343, b => 344, p => False), (a => 345, b => 346, p => False), (a => 347, b => 348, p => False), (a => 349, b => 350, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 258, p => True ), (a => 2  , b => 257, p => True ), (a => 3  , b => 256, p => True ), (a => 124, b => 255, p => True ), (a => 125, b => 128, p => True ), (a => 126, b => 127, p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 26 , b => 28 , p => False), (a => 30 , b => 32 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 42 , b => 44 , p => False), (a => 46 , b => 48 , p => False), (a => 50 , b => 52 , p => False), (a => 54 , b => 56 , p => False), (a => 58 , b => 60 , p => False), (a => 62 , b => 64 , p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 74 , b => 76 , p => False), (a => 78 , b => 80 , p => False), (a => 82 , b => 84 , p => False), (a => 86 , b => 88 , p => False), (a => 90 , b => 92 , p => False), (a => 94 , b => 96 , p => False), (a => 98 , b => 100, p => False), (a => 102, b => 104, p => False), (a => 106, b => 108, p => False), (a => 110, b => 112, p => False), (a => 114, b => 116, p => False), (a => 118, b => 120, p => False), (a => 122, b => 124, p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 27 , b => 29 , p => False), (a => 31 , b => 33 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 43 , b => 45 , p => False), (a => 47 , b => 49 , p => False), (a => 51 , b => 53 , p => False), (a => 55 , b => 57 , p => False), (a => 59 , b => 61 , p => False), (a => 63 , b => 65 , p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 75 , b => 77 , p => False), (a => 79 , b => 81 , p => False), (a => 83 , b => 85 , p => False), (a => 87 , b => 89 , p => False), (a => 91 , b => 93 , p => False), (a => 95 , b => 97 , p => False), (a => 99 , b => 101, p => False), (a => 103, b => 105, p => False), (a => 107, b => 109, p => False), (a => 111, b => 113, p => False), (a => 115, b => 117, p => False), (a => 119, b => 121, p => False), (a => 123, b => 125, p => False), (a => 288, b => 320, p => False), (a => 304, b => 336, p => False), (a => 296, b => 328, p => False), (a => 312, b => 344, p => False), (a => 292, b => 324, p => False), (a => 308, b => 340, p => False), (a => 300, b => 332, p => False), (a => 316, b => 348, p => False), (a => 290, b => 322, p => False), (a => 306, b => 338, p => False), (a => 298, b => 330, p => False), (a => 314, b => 346, p => False), (a => 294, b => 326, p => False), (a => 310, b => 342, p => False), (a => 302, b => 334, p => False), (a => 318, b => 350, p => False), (a => 289, b => 321, p => False), (a => 305, b => 337, p => False), (a => 297, b => 329, p => False), (a => 313, b => 345, p => False), (a => 293, b => 325, p => False), (a => 309, b => 341, p => False), (a => 301, b => 333, p => False), (a => 317, b => 349, p => False), (a => 291, b => 323, p => False), (a => 307, b => 339, p => False), (a => 299, b => 331, p => False), (a => 315, b => 347, p => False), (a => 295, b => 327, p => False), (a => 311, b => 343, p => False), (a => 303, b => 335, p => False), (a => 319, b => 351, p => False), (a => 0  , b => 287, p => True ), (a => 1  , b => 286, p => True ), (a => 126, b => 285, p => True ), (a => 127, b => 284, p => True ), (a => 128, b => 283, p => True ), (a => 129, b => 282, p => True ), (a => 130, b => 281, p => True ), (a => 131, b => 280, p => True ), (a => 132, b => 279, p => True ), (a => 133, b => 278, p => True ), (a => 134, b => 277, p => True ), (a => 135, b => 276, p => True ), (a => 136, b => 275, p => True ), (a => 137, b => 274, p => True ), (a => 138, b => 273, p => True ), (a => 139, b => 272, p => True ), (a => 140, b => 271, p => True ), (a => 141, b => 270, p => True ), (a => 142, b => 269, p => True ), (a => 143, b => 268, p => True ), (a => 144, b => 267, p => True ), (a => 145, b => 266, p => True ), (a => 146, b => 265, p => True ), (a => 147, b => 264, p => True ), (a => 148, b => 263, p => True ), (a => 149, b => 262, p => True ), (a => 150, b => 261, p => True ), (a => 151, b => 260, p => True ), (a => 152, b => 259, p => True ), (a => 153, b => 258, p => True ), (a => 154, b => 257, p => True ), (a => 155, b => 256, p => True ), (a => 156, b => 255, p => True ), (a => 157, b => 254, p => True ), (a => 158, b => 253, p => True ), (a => 159, b => 252, p => True ), (a => 160, b => 251, p => True ), (a => 161, b => 250, p => True ), (a => 162, b => 249, p => True ), (a => 163, b => 248, p => True ), (a => 164, b => 247, p => True ), (a => 165, b => 246, p => True ), (a => 166, b => 245, p => True ), (a => 167, b => 244, p => True ), (a => 168, b => 243, p => True ), (a => 169, b => 242, p => True ), (a => 170, b => 241, p => True ), (a => 171, b => 240, p => True ), (a => 172, b => 239, p => True ), (a => 173, b => 238, p => True ), (a => 174, b => 237, p => True ), (a => 175, b => 236, p => True ), (a => 176, b => 235, p => True ), (a => 177, b => 234, p => True ), (a => 178, b => 233, p => True ), (a => 179, b => 232, p => True ), (a => 180, b => 231, p => True ), (a => 181, b => 230, p => True ), (a => 182, b => 229, p => True ), (a => 183, b => 228, p => True ), (a => 184, b => 227, p => True ), (a => 185, b => 226, p => True ), (a => 186, b => 225, p => True ), (a => 187, b => 224, p => True ), (a => 188, b => 223, p => True ), (a => 189, b => 222, p => True ), (a => 190, b => 221, p => True ), (a => 191, b => 220, p => True ), (a => 192, b => 219, p => True ), (a => 193, b => 218, p => True ), (a => 194, b => 217, p => True ), (a => 195, b => 216, p => True ), (a => 196, b => 215, p => True ), (a => 197, b => 214, p => True ), (a => 198, b => 213, p => True ), (a => 199, b => 212, p => True ), (a => 200, b => 211, p => True ), (a => 201, b => 210, p => True ), (a => 202, b => 209, p => True ), (a => 203, b => 208, p => True ), (a => 204, b => 207, p => True ), (a => 205, b => 206, p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 25 , b => 26 , p => False), (a => 27 , b => 28 , p => False), (a => 29 , b => 30 , p => False), (a => 31 , b => 32 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 41 , b => 42 , p => False), (a => 43 , b => 44 , p => False), (a => 45 , b => 46 , p => False), (a => 47 , b => 48 , p => False), (a => 49 , b => 50 , p => False), (a => 51 , b => 52 , p => False), (a => 53 , b => 54 , p => False), (a => 55 , b => 56 , p => False), (a => 57 , b => 58 , p => False), (a => 59 , b => 60 , p => False), (a => 61 , b => 62 , p => False), (a => 63 , b => 64 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 73 , b => 74 , p => False), (a => 75 , b => 76 , p => False), (a => 77 , b => 78 , p => False), (a => 79 , b => 80 , p => False), (a => 81 , b => 82 , p => False), (a => 83 , b => 84 , p => False), (a => 85 , b => 86 , p => False), (a => 87 , b => 88 , p => False), (a => 89 , b => 90 , p => False), (a => 91 , b => 92 , p => False), (a => 93 , b => 94 , p => False), (a => 95 , b => 96 , p => False), (a => 97 , b => 98 , p => False), (a => 99 , b => 100, p => False), (a => 101, b => 102, p => False), (a => 103, b => 104, p => False), (a => 105, b => 106, p => False), (a => 107, b => 108, p => False), (a => 109, b => 110, p => False), (a => 111, b => 112, p => False), (a => 113, b => 114, p => False), (a => 115, b => 116, p => False), (a => 117, b => 118, p => False), (a => 119, b => 120, p => False), (a => 121, b => 122, p => False), (a => 123, b => 124, p => False), (a => 125, b => 126, p => False), (a => 272, b => 288, p => False), (a => 304, b => 320, p => False), (a => 280, b => 296, p => False), (a => 312, b => 328, p => False), (a => 276, b => 292, p => False), (a => 308, b => 324, p => False), (a => 284, b => 300, p => False), (a => 316, b => 332, p => False), (a => 274, b => 290, p => False), (a => 306, b => 322, p => False), (a => 282, b => 298, p => False), (a => 314, b => 330, p => False), (a => 278, b => 294, p => False), (a => 310, b => 326, p => False), (a => 286, b => 302, p => False), (a => 318, b => 334, p => False), (a => 273, b => 289, p => False), (a => 305, b => 321, p => False), (a => 281, b => 297, p => False), (a => 313, b => 329, p => False), (a => 277, b => 293, p => False), (a => 309, b => 325, p => False), (a => 285, b => 301, p => False), (a => 317, b => 333, p => False), (a => 275, b => 291, p => False), (a => 307, b => 323, p => False), (a => 283, b => 299, p => False), (a => 315, b => 331, p => False), (a => 279, b => 295, p => False), (a => 311, b => 327, p => False), (a => 287, b => 303, p => False), (a => 319, b => 335, p => False), (a => 0  , b => 351, p => True ), (a => 127, b => 350, p => True ), (a => 128, b => 349, p => True ), (a => 129, b => 348, p => True ), (a => 130, b => 347, p => True ), (a => 131, b => 346, p => True ), (a => 132, b => 345, p => True ), (a => 133, b => 344, p => True ), (a => 134, b => 343, p => True ), (a => 135, b => 342, p => True ), (a => 136, b => 341, p => True ), (a => 137, b => 340, p => True ), (a => 138, b => 339, p => True ), (a => 139, b => 338, p => True ), (a => 140, b => 337, p => True ), (a => 141, b => 336, p => True ), (a => 142, b => 271, p => True ), (a => 143, b => 270, p => True ), (a => 144, b => 269, p => True ), (a => 145, b => 268, p => True ), (a => 146, b => 267, p => True ), (a => 147, b => 266, p => True ), (a => 148, b => 265, p => True ), (a => 149, b => 264, p => True ), (a => 150, b => 263, p => True ), (a => 151, b => 262, p => True ), (a => 152, b => 261, p => True ), (a => 153, b => 260, p => True ), (a => 154, b => 259, p => True ), (a => 155, b => 258, p => True ), (a => 156, b => 257, p => True ), (a => 157, b => 256, p => True ), (a => 158, b => 255, p => True ), (a => 159, b => 254, p => True ), (a => 160, b => 253, p => True ), (a => 161, b => 252, p => True ), (a => 162, b => 251, p => True ), (a => 163, b => 250, p => True ), (a => 164, b => 249, p => True ), (a => 165, b => 248, p => True ), (a => 166, b => 247, p => True ), (a => 167, b => 246, p => True ), (a => 168, b => 245, p => True ), (a => 169, b => 244, p => True ), (a => 170, b => 243, p => True ), (a => 171, b => 242, p => True ), (a => 172, b => 241, p => True ), (a => 173, b => 240, p => True ), (a => 174, b => 239, p => True ), (a => 175, b => 238, p => True ), (a => 176, b => 237, p => True ), (a => 177, b => 236, p => True ), (a => 178, b => 235, p => True ), (a => 179, b => 234, p => True ), (a => 180, b => 233, p => True ), (a => 181, b => 232, p => True ), (a => 182, b => 231, p => True ), (a => 183, b => 230, p => True ), (a => 184, b => 229, p => True ), (a => 185, b => 228, p => True ), (a => 186, b => 227, p => True ), (a => 187, b => 226, p => True ), (a => 188, b => 225, p => True ), (a => 189, b => 224, p => True ), (a => 190, b => 223, p => True ), (a => 191, b => 222, p => True ), (a => 192, b => 221, p => True ), (a => 193, b => 220, p => True ), (a => 194, b => 219, p => True ), (a => 195, b => 218, p => True ), (a => 196, b => 217, p => True ), (a => 197, b => 216, p => True ), (a => 198, b => 215, p => True ), (a => 199, b => 214, p => True ), (a => 200, b => 213, p => True ), (a => 201, b => 212, p => True ), (a => 202, b => 211, p => True ), (a => 203, b => 210, p => True ), (a => 204, b => 209, p => True ), (a => 205, b => 208, p => True ), (a => 206, b => 207, p => True )),
                    ((a => 64 , b => 192, p => False), (a => 32 , b => 160, p => False), (a => 96 , b => 224, p => False), (a => 16 , b => 144, p => False), (a => 80 , b => 208, p => False), (a => 48 , b => 176, p => False), (a => 112, b => 240, p => False), (a => 8  , b => 136, p => False), (a => 72 , b => 200, p => False), (a => 40 , b => 168, p => False), (a => 104, b => 232, p => False), (a => 24 , b => 152, p => False), (a => 88 , b => 216, p => False), (a => 56 , b => 184, p => False), (a => 120, b => 248, p => False), (a => 4  , b => 132, p => False), (a => 68 , b => 196, p => False), (a => 36 , b => 164, p => False), (a => 100, b => 228, p => False), (a => 20 , b => 148, p => False), (a => 84 , b => 212, p => False), (a => 52 , b => 180, p => False), (a => 116, b => 244, p => False), (a => 12 , b => 140, p => False), (a => 76 , b => 204, p => False), (a => 44 , b => 172, p => False), (a => 108, b => 236, p => False), (a => 28 , b => 156, p => False), (a => 92 , b => 220, p => False), (a => 60 , b => 188, p => False), (a => 124, b => 252, p => False), (a => 2  , b => 130, p => False), (a => 66 , b => 194, p => False), (a => 34 , b => 162, p => False), (a => 98 , b => 226, p => False), (a => 18 , b => 146, p => False), (a => 82 , b => 210, p => False), (a => 50 , b => 178, p => False), (a => 114, b => 242, p => False), (a => 10 , b => 138, p => False), (a => 74 , b => 202, p => False), (a => 42 , b => 170, p => False), (a => 106, b => 234, p => False), (a => 26 , b => 154, p => False), (a => 90 , b => 218, p => False), (a => 58 , b => 186, p => False), (a => 122, b => 250, p => False), (a => 6  , b => 134, p => False), (a => 70 , b => 198, p => False), (a => 38 , b => 166, p => False), (a => 102, b => 230, p => False), (a => 22 , b => 150, p => False), (a => 86 , b => 214, p => False), (a => 54 , b => 182, p => False), (a => 118, b => 246, p => False), (a => 14 , b => 142, p => False), (a => 78 , b => 206, p => False), (a => 46 , b => 174, p => False), (a => 110, b => 238, p => False), (a => 30 , b => 158, p => False), (a => 94 , b => 222, p => False), (a => 62 , b => 190, p => False), (a => 126, b => 254, p => False), (a => 1  , b => 129, p => False), (a => 65 , b => 193, p => False), (a => 33 , b => 161, p => False), (a => 97 , b => 225, p => False), (a => 17 , b => 145, p => False), (a => 81 , b => 209, p => False), (a => 49 , b => 177, p => False), (a => 113, b => 241, p => False), (a => 9  , b => 137, p => False), (a => 73 , b => 201, p => False), (a => 41 , b => 169, p => False), (a => 105, b => 233, p => False), (a => 25 , b => 153, p => False), (a => 89 , b => 217, p => False), (a => 57 , b => 185, p => False), (a => 121, b => 249, p => False), (a => 5  , b => 133, p => False), (a => 69 , b => 197, p => False), (a => 37 , b => 165, p => False), (a => 101, b => 229, p => False), (a => 21 , b => 149, p => False), (a => 85 , b => 213, p => False), (a => 53 , b => 181, p => False), (a => 117, b => 245, p => False), (a => 13 , b => 141, p => False), (a => 77 , b => 205, p => False), (a => 45 , b => 173, p => False), (a => 109, b => 237, p => False), (a => 29 , b => 157, p => False), (a => 93 , b => 221, p => False), (a => 61 , b => 189, p => False), (a => 125, b => 253, p => False), (a => 3  , b => 131, p => False), (a => 67 , b => 195, p => False), (a => 35 , b => 163, p => False), (a => 99 , b => 227, p => False), (a => 19 , b => 147, p => False), (a => 83 , b => 211, p => False), (a => 51 , b => 179, p => False), (a => 115, b => 243, p => False), (a => 11 , b => 139, p => False), (a => 75 , b => 203, p => False), (a => 43 , b => 171, p => False), (a => 107, b => 235, p => False), (a => 27 , b => 155, p => False), (a => 91 , b => 219, p => False), (a => 59 , b => 187, p => False), (a => 123, b => 251, p => False), (a => 7  , b => 135, p => False), (a => 71 , b => 199, p => False), (a => 39 , b => 167, p => False), (a => 103, b => 231, p => False), (a => 23 , b => 151, p => False), (a => 87 , b => 215, p => False), (a => 55 , b => 183, p => False), (a => 119, b => 247, p => False), (a => 15 , b => 143, p => False), (a => 79 , b => 207, p => False), (a => 47 , b => 175, p => False), (a => 111, b => 239, p => False), (a => 31 , b => 159, p => False), (a => 95 , b => 223, p => False), (a => 63 , b => 191, p => False), (a => 264, b => 272, p => False), (a => 280, b => 288, p => False), (a => 296, b => 304, p => False), (a => 312, b => 320, p => False), (a => 328, b => 336, p => False), (a => 268, b => 276, p => False), (a => 284, b => 292, p => False), (a => 316, b => 324, p => False), (a => 266, b => 274, p => False), (a => 282, b => 290, p => False), (a => 298, b => 306, p => False), (a => 314, b => 322, p => False), (a => 330, b => 338, p => False), (a => 270, b => 278, p => False), (a => 286, b => 294, p => False), (a => 318, b => 326, p => False), (a => 265, b => 273, p => False), (a => 281, b => 289, p => False), (a => 297, b => 305, p => False), (a => 313, b => 321, p => False), (a => 329, b => 337, p => False), (a => 269, b => 277, p => False), (a => 285, b => 293, p => False), (a => 317, b => 325, p => False), (a => 267, b => 275, p => False), (a => 283, b => 291, p => False), (a => 299, b => 307, p => False), (a => 315, b => 323, p => False), (a => 331, b => 339, p => False), (a => 271, b => 279, p => False), (a => 287, b => 295, p => False), (a => 319, b => 327, p => False), (a => 0  , b => 351, p => True ), (a => 127, b => 350, p => True ), (a => 128, b => 349, p => True ), (a => 255, b => 348, p => True ), (a => 256, b => 347, p => True ), (a => 257, b => 346, p => True ), (a => 258, b => 345, p => True ), (a => 259, b => 344, p => True ), (a => 260, b => 343, p => True ), (a => 261, b => 342, p => True ), (a => 262, b => 341, p => True ), (a => 263, b => 340, p => True ), (a => 300, b => 335, p => True ), (a => 301, b => 334, p => True ), (a => 302, b => 333, p => True ), (a => 303, b => 332, p => True ), (a => 308, b => 311, p => True ), (a => 309, b => 310, p => True )),
                    ((a => 64 , b => 128, p => False), (a => 96 , b => 160, p => False), (a => 80 , b => 144, p => False), (a => 112, b => 176, p => False), (a => 72 , b => 136, p => False), (a => 104, b => 168, p => False), (a => 88 , b => 152, p => False), (a => 120, b => 184, p => False), (a => 68 , b => 132, p => False), (a => 100, b => 164, p => False), (a => 84 , b => 148, p => False), (a => 116, b => 180, p => False), (a => 76 , b => 140, p => False), (a => 108, b => 172, p => False), (a => 92 , b => 156, p => False), (a => 124, b => 188, p => False), (a => 66 , b => 130, p => False), (a => 98 , b => 162, p => False), (a => 82 , b => 146, p => False), (a => 114, b => 178, p => False), (a => 74 , b => 138, p => False), (a => 106, b => 170, p => False), (a => 90 , b => 154, p => False), (a => 122, b => 186, p => False), (a => 70 , b => 134, p => False), (a => 102, b => 166, p => False), (a => 86 , b => 150, p => False), (a => 118, b => 182, p => False), (a => 78 , b => 142, p => False), (a => 110, b => 174, p => False), (a => 94 , b => 158, p => False), (a => 126, b => 190, p => False), (a => 65 , b => 129, p => False), (a => 97 , b => 161, p => False), (a => 81 , b => 145, p => False), (a => 113, b => 177, p => False), (a => 73 , b => 137, p => False), (a => 105, b => 169, p => False), (a => 89 , b => 153, p => False), (a => 121, b => 185, p => False), (a => 69 , b => 133, p => False), (a => 101, b => 165, p => False), (a => 85 , b => 149, p => False), (a => 117, b => 181, p => False), (a => 77 , b => 141, p => False), (a => 109, b => 173, p => False), (a => 93 , b => 157, p => False), (a => 125, b => 189, p => False), (a => 67 , b => 131, p => False), (a => 99 , b => 163, p => False), (a => 83 , b => 147, p => False), (a => 115, b => 179, p => False), (a => 75 , b => 139, p => False), (a => 107, b => 171, p => False), (a => 91 , b => 155, p => False), (a => 123, b => 187, p => False), (a => 71 , b => 135, p => False), (a => 103, b => 167, p => False), (a => 87 , b => 151, p => False), (a => 119, b => 183, p => False), (a => 79 , b => 143, p => False), (a => 111, b => 175, p => False), (a => 95 , b => 159, p => False), (a => 127, b => 191, p => False), (a => 260, b => 264, p => False), (a => 268, b => 272, p => False), (a => 276, b => 280, p => False), (a => 284, b => 288, p => False), (a => 292, b => 296, p => False), (a => 316, b => 320, p => False), (a => 324, b => 328, p => False), (a => 262, b => 266, p => False), (a => 270, b => 274, p => False), (a => 278, b => 282, p => False), (a => 286, b => 290, p => False), (a => 294, b => 298, p => False), (a => 318, b => 322, p => False), (a => 326, b => 330, p => False), (a => 261, b => 265, p => False), (a => 269, b => 273, p => False), (a => 277, b => 281, p => False), (a => 285, b => 289, p => False), (a => 293, b => 297, p => False), (a => 317, b => 321, p => False), (a => 325, b => 329, p => False), (a => 263, b => 267, p => False), (a => 271, b => 275, p => False), (a => 279, b => 283, p => False), (a => 287, b => 291, p => False), (a => 295, b => 299, p => False), (a => 319, b => 323, p => False), (a => 327, b => 331, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 343, p => True ), (a => 9  , b => 342, p => True ), (a => 10 , b => 341, p => True ), (a => 11 , b => 340, p => True ), (a => 12 , b => 339, p => True ), (a => 13 , b => 338, p => True ), (a => 14 , b => 337, p => True ), (a => 15 , b => 336, p => True ), (a => 16 , b => 335, p => True ), (a => 17 , b => 334, p => True ), (a => 18 , b => 333, p => True ), (a => 19 , b => 332, p => True ), (a => 20 , b => 315, p => True ), (a => 21 , b => 314, p => True ), (a => 22 , b => 313, p => True ), (a => 23 , b => 312, p => True ), (a => 24 , b => 311, p => True ), (a => 25 , b => 310, p => True ), (a => 26 , b => 309, p => True ), (a => 27 , b => 308, p => True ), (a => 28 , b => 307, p => True ), (a => 29 , b => 306, p => True ), (a => 30 , b => 305, p => True ), (a => 31 , b => 304, p => True ), (a => 32 , b => 303, p => True ), (a => 33 , b => 302, p => True ), (a => 34 , b => 301, p => True ), (a => 35 , b => 300, p => True ), (a => 36 , b => 259, p => True ), (a => 37 , b => 258, p => True ), (a => 38 , b => 257, p => True ), (a => 39 , b => 256, p => True ), (a => 40 , b => 255, p => True ), (a => 41 , b => 254, p => True ), (a => 42 , b => 253, p => True ), (a => 43 , b => 252, p => True ), (a => 44 , b => 251, p => True ), (a => 45 , b => 250, p => True ), (a => 46 , b => 249, p => True ), (a => 47 , b => 248, p => True ), (a => 48 , b => 247, p => True ), (a => 49 , b => 246, p => True ), (a => 50 , b => 245, p => True ), (a => 51 , b => 244, p => True ), (a => 52 , b => 243, p => True ), (a => 53 , b => 242, p => True ), (a => 54 , b => 241, p => True ), (a => 55 , b => 240, p => True ), (a => 56 , b => 239, p => True ), (a => 57 , b => 238, p => True ), (a => 58 , b => 237, p => True ), (a => 59 , b => 236, p => True ), (a => 60 , b => 235, p => True ), (a => 61 , b => 234, p => True ), (a => 62 , b => 233, p => True ), (a => 63 , b => 232, p => True ), (a => 192, b => 231, p => True ), (a => 193, b => 230, p => True ), (a => 194, b => 229, p => True ), (a => 195, b => 228, p => True ), (a => 196, b => 227, p => True ), (a => 197, b => 226, p => True ), (a => 198, b => 225, p => True ), (a => 199, b => 224, p => True ), (a => 200, b => 223, p => True ), (a => 201, b => 222, p => True ), (a => 202, b => 221, p => True ), (a => 203, b => 220, p => True ), (a => 204, b => 219, p => True ), (a => 205, b => 218, p => True ), (a => 206, b => 217, p => True ), (a => 207, b => 216, p => True ), (a => 208, b => 215, p => True ), (a => 209, b => 214, p => True ), (a => 210, b => 213, p => True ), (a => 211, b => 212, p => True )),
                    ((a => 32 , b => 64 , p => False), (a => 96 , b => 128, p => False), (a => 160, b => 192, p => False), (a => 48 , b => 80 , p => False), (a => 112, b => 144, p => False), (a => 40 , b => 72 , p => False), (a => 104, b => 136, p => False), (a => 56 , b => 88 , p => False), (a => 120, b => 152, p => False), (a => 36 , b => 68 , p => False), (a => 100, b => 132, p => False), (a => 52 , b => 84 , p => False), (a => 116, b => 148, p => False), (a => 44 , b => 76 , p => False), (a => 108, b => 140, p => False), (a => 60 , b => 92 , p => False), (a => 124, b => 156, p => False), (a => 34 , b => 66 , p => False), (a => 98 , b => 130, p => False), (a => 162, b => 194, p => False), (a => 50 , b => 82 , p => False), (a => 114, b => 146, p => False), (a => 42 , b => 74 , p => False), (a => 106, b => 138, p => False), (a => 58 , b => 90 , p => False), (a => 122, b => 154, p => False), (a => 38 , b => 70 , p => False), (a => 102, b => 134, p => False), (a => 54 , b => 86 , p => False), (a => 118, b => 150, p => False), (a => 46 , b => 78 , p => False), (a => 110, b => 142, p => False), (a => 62 , b => 94 , p => False), (a => 126, b => 158, p => False), (a => 33 , b => 65 , p => False), (a => 97 , b => 129, p => False), (a => 161, b => 193, p => False), (a => 49 , b => 81 , p => False), (a => 113, b => 145, p => False), (a => 41 , b => 73 , p => False), (a => 105, b => 137, p => False), (a => 57 , b => 89 , p => False), (a => 121, b => 153, p => False), (a => 37 , b => 69 , p => False), (a => 101, b => 133, p => False), (a => 53 , b => 85 , p => False), (a => 117, b => 149, p => False), (a => 45 , b => 77 , p => False), (a => 109, b => 141, p => False), (a => 61 , b => 93 , p => False), (a => 125, b => 157, p => False), (a => 35 , b => 67 , p => False), (a => 99 , b => 131, p => False), (a => 163, b => 195, p => False), (a => 51 , b => 83 , p => False), (a => 115, b => 147, p => False), (a => 43 , b => 75 , p => False), (a => 107, b => 139, p => False), (a => 59 , b => 91 , p => False), (a => 123, b => 155, p => False), (a => 39 , b => 71 , p => False), (a => 103, b => 135, p => False), (a => 55 , b => 87 , p => False), (a => 119, b => 151, p => False), (a => 47 , b => 79 , p => False), (a => 111, b => 143, p => False), (a => 63 , b => 95 , p => False), (a => 127, b => 159, p => False), (a => 258, b => 260, p => False), (a => 262, b => 264, p => False), (a => 266, b => 268, p => False), (a => 270, b => 272, p => False), (a => 274, b => 276, p => False), (a => 278, b => 280, p => False), (a => 286, b => 288, p => False), (a => 290, b => 292, p => False), (a => 294, b => 296, p => False), (a => 318, b => 320, p => False), (a => 322, b => 324, p => False), (a => 326, b => 328, p => False), (a => 259, b => 261, p => False), (a => 263, b => 265, p => False), (a => 267, b => 269, p => False), (a => 271, b => 273, p => False), (a => 275, b => 277, p => False), (a => 279, b => 281, p => False), (a => 287, b => 289, p => False), (a => 291, b => 293, p => False), (a => 295, b => 297, p => False), (a => 319, b => 321, p => False), (a => 323, b => 325, p => False), (a => 327, b => 329, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 343, p => True ), (a => 9  , b => 342, p => True ), (a => 10 , b => 341, p => True ), (a => 11 , b => 340, p => True ), (a => 12 , b => 339, p => True ), (a => 13 , b => 338, p => True ), (a => 14 , b => 337, p => True ), (a => 15 , b => 336, p => True ), (a => 16 , b => 335, p => True ), (a => 17 , b => 334, p => True ), (a => 18 , b => 333, p => True ), (a => 19 , b => 332, p => True ), (a => 20 , b => 331, p => True ), (a => 21 , b => 330, p => True ), (a => 22 , b => 317, p => True ), (a => 23 , b => 316, p => True ), (a => 24 , b => 315, p => True ), (a => 25 , b => 314, p => True ), (a => 26 , b => 313, p => True ), (a => 27 , b => 312, p => True ), (a => 28 , b => 311, p => True ), (a => 29 , b => 310, p => True ), (a => 30 , b => 309, p => True ), (a => 31 , b => 308, p => True ), (a => 164, b => 307, p => True ), (a => 165, b => 306, p => True ), (a => 166, b => 305, p => True ), (a => 167, b => 304, p => True ), (a => 168, b => 303, p => True ), (a => 169, b => 302, p => True ), (a => 170, b => 301, p => True ), (a => 171, b => 300, p => True ), (a => 172, b => 299, p => True ), (a => 173, b => 298, p => True ), (a => 174, b => 285, p => True ), (a => 175, b => 284, p => True ), (a => 176, b => 283, p => True ), (a => 177, b => 282, p => True ), (a => 178, b => 257, p => True ), (a => 179, b => 256, p => True ), (a => 180, b => 255, p => True ), (a => 181, b => 254, p => True ), (a => 182, b => 253, p => True ), (a => 183, b => 252, p => True ), (a => 184, b => 251, p => True ), (a => 185, b => 250, p => True ), (a => 186, b => 249, p => True ), (a => 187, b => 248, p => True ), (a => 188, b => 247, p => True ), (a => 189, b => 246, p => True ), (a => 190, b => 245, p => True ), (a => 191, b => 244, p => True ), (a => 196, b => 243, p => True ), (a => 197, b => 242, p => True ), (a => 198, b => 241, p => True ), (a => 199, b => 240, p => True ), (a => 200, b => 239, p => True ), (a => 201, b => 238, p => True ), (a => 202, b => 237, p => True ), (a => 203, b => 236, p => True ), (a => 204, b => 235, p => True ), (a => 205, b => 234, p => True ), (a => 206, b => 233, p => True ), (a => 207, b => 232, p => True ), (a => 208, b => 231, p => True ), (a => 209, b => 230, p => True ), (a => 210, b => 229, p => True ), (a => 211, b => 228, p => True ), (a => 212, b => 227, p => True ), (a => 213, b => 226, p => True ), (a => 214, b => 225, p => True ), (a => 215, b => 224, p => True ), (a => 216, b => 223, p => True ), (a => 217, b => 222, p => True ), (a => 218, b => 221, p => True ), (a => 219, b => 220, p => True )),
                    ((a => 16 , b => 32 , p => False), (a => 48 , b => 64 , p => False), (a => 80 , b => 96 , p => False), (a => 112, b => 128, p => False), (a => 144, b => 160, p => False), (a => 24 , b => 40 , p => False), (a => 56 , b => 72 , p => False), (a => 120, b => 136, p => False), (a => 20 , b => 36 , p => False), (a => 52 , b => 68 , p => False), (a => 116, b => 132, p => False), (a => 28 , b => 44 , p => False), (a => 60 , b => 76 , p => False), (a => 124, b => 140, p => False), (a => 18 , b => 34 , p => False), (a => 50 , b => 66 , p => False), (a => 82 , b => 98 , p => False), (a => 114, b => 130, p => False), (a => 146, b => 162, p => False), (a => 26 , b => 42 , p => False), (a => 58 , b => 74 , p => False), (a => 122, b => 138, p => False), (a => 22 , b => 38 , p => False), (a => 54 , b => 70 , p => False), (a => 118, b => 134, p => False), (a => 30 , b => 46 , p => False), (a => 62 , b => 78 , p => False), (a => 126, b => 142, p => False), (a => 17 , b => 33 , p => False), (a => 49 , b => 65 , p => False), (a => 81 , b => 97 , p => False), (a => 113, b => 129, p => False), (a => 145, b => 161, p => False), (a => 25 , b => 41 , p => False), (a => 57 , b => 73 , p => False), (a => 121, b => 137, p => False), (a => 21 , b => 37 , p => False), (a => 53 , b => 69 , p => False), (a => 117, b => 133, p => False), (a => 29 , b => 45 , p => False), (a => 61 , b => 77 , p => False), (a => 125, b => 141, p => False), (a => 19 , b => 35 , p => False), (a => 51 , b => 67 , p => False), (a => 83 , b => 99 , p => False), (a => 115, b => 131, p => False), (a => 147, b => 163, p => False), (a => 27 , b => 43 , p => False), (a => 59 , b => 75 , p => False), (a => 123, b => 139, p => False), (a => 23 , b => 39 , p => False), (a => 55 , b => 71 , p => False), (a => 119, b => 135, p => False), (a => 31 , b => 47 , p => False), (a => 63 , b => 79 , p => False), (a => 127, b => 143, p => False), (a => 257, b => 258, p => False), (a => 259, b => 260, p => False), (a => 261, b => 262, p => False), (a => 263, b => 264, p => False), (a => 265, b => 266, p => False), (a => 267, b => 268, p => False), (a => 269, b => 270, p => False), (a => 271, b => 272, p => False), (a => 273, b => 274, p => False), (a => 275, b => 276, p => False), (a => 277, b => 278, p => False), (a => 279, b => 280, p => False), (a => 287, b => 288, p => False), (a => 289, b => 290, p => False), (a => 291, b => 292, p => False), (a => 293, b => 294, p => False), (a => 295, b => 296, p => False), (a => 319, b => 320, p => False), (a => 321, b => 322, p => False), (a => 323, b => 324, p => False), (a => 325, b => 326, p => False), (a => 327, b => 328, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 343, p => True ), (a => 9  , b => 342, p => True ), (a => 10 , b => 341, p => True ), (a => 11 , b => 340, p => True ), (a => 12 , b => 339, p => True ), (a => 13 , b => 338, p => True ), (a => 14 , b => 337, p => True ), (a => 15 , b => 336, p => True ), (a => 84 , b => 335, p => True ), (a => 85 , b => 334, p => True ), (a => 86 , b => 333, p => True ), (a => 87 , b => 332, p => True ), (a => 88 , b => 331, p => True ), (a => 89 , b => 330, p => True ), (a => 90 , b => 329, p => True ), (a => 91 , b => 318, p => True ), (a => 92 , b => 317, p => True ), (a => 93 , b => 316, p => True ), (a => 94 , b => 315, p => True ), (a => 95 , b => 314, p => True ), (a => 100, b => 313, p => True ), (a => 101, b => 312, p => True ), (a => 102, b => 311, p => True ), (a => 103, b => 310, p => True ), (a => 104, b => 309, p => True ), (a => 105, b => 308, p => True ), (a => 106, b => 307, p => True ), (a => 107, b => 306, p => True ), (a => 108, b => 305, p => True ), (a => 109, b => 304, p => True ), (a => 110, b => 303, p => True ), (a => 111, b => 302, p => True ), (a => 148, b => 301, p => True ), (a => 149, b => 300, p => True ), (a => 150, b => 299, p => True ), (a => 151, b => 298, p => True ), (a => 152, b => 297, p => True ), (a => 153, b => 286, p => True ), (a => 154, b => 285, p => True ), (a => 155, b => 284, p => True ), (a => 156, b => 283, p => True ), (a => 157, b => 282, p => True ), (a => 158, b => 281, p => True ), (a => 159, b => 256, p => True ), (a => 164, b => 255, p => True ), (a => 165, b => 254, p => True ), (a => 166, b => 253, p => True ), (a => 167, b => 252, p => True ), (a => 168, b => 251, p => True ), (a => 169, b => 250, p => True ), (a => 170, b => 249, p => True ), (a => 171, b => 248, p => True ), (a => 172, b => 247, p => True ), (a => 173, b => 246, p => True ), (a => 174, b => 245, p => True ), (a => 175, b => 244, p => True ), (a => 176, b => 243, p => True ), (a => 177, b => 242, p => True ), (a => 178, b => 241, p => True ), (a => 179, b => 240, p => True ), (a => 180, b => 239, p => True ), (a => 181, b => 238, p => True ), (a => 182, b => 237, p => True ), (a => 183, b => 236, p => True ), (a => 184, b => 235, p => True ), (a => 185, b => 234, p => True ), (a => 186, b => 233, p => True ), (a => 187, b => 232, p => True ), (a => 188, b => 231, p => True ), (a => 189, b => 230, p => True ), (a => 190, b => 229, p => True ), (a => 191, b => 228, p => True ), (a => 192, b => 227, p => True ), (a => 193, b => 226, p => True ), (a => 194, b => 225, p => True ), (a => 195, b => 224, p => True ), (a => 196, b => 223, p => True ), (a => 197, b => 222, p => True ), (a => 198, b => 221, p => True ), (a => 199, b => 220, p => True ), (a => 200, b => 219, p => True ), (a => 201, b => 218, p => True ), (a => 202, b => 217, p => True ), (a => 203, b => 216, p => True ), (a => 204, b => 215, p => True ), (a => 205, b => 214, p => True ), (a => 206, b => 213, p => True ), (a => 207, b => 212, p => True ), (a => 208, b => 211, p => True ), (a => 209, b => 210, p => True )),
                    ((a => 8  , b => 16 , p => False), (a => 24 , b => 32 , p => False), (a => 40 , b => 48 , p => False), (a => 56 , b => 64 , p => False), (a => 72 , b => 80 , p => False), (a => 120, b => 128, p => False), (a => 136, b => 144, p => False), (a => 12 , b => 20 , p => False), (a => 28 , b => 36 , p => False), (a => 60 , b => 68 , p => False), (a => 124, b => 132, p => False), (a => 10 , b => 18 , p => False), (a => 26 , b => 34 , p => False), (a => 42 , b => 50 , p => False), (a => 58 , b => 66 , p => False), (a => 74 , b => 82 , p => False), (a => 122, b => 130, p => False), (a => 138, b => 146, p => False), (a => 14 , b => 22 , p => False), (a => 30 , b => 38 , p => False), (a => 62 , b => 70 , p => False), (a => 126, b => 134, p => False), (a => 9  , b => 17 , p => False), (a => 25 , b => 33 , p => False), (a => 41 , b => 49 , p => False), (a => 57 , b => 65 , p => False), (a => 73 , b => 81 , p => False), (a => 121, b => 129, p => False), (a => 137, b => 145, p => False), (a => 13 , b => 21 , p => False), (a => 29 , b => 37 , p => False), (a => 61 , b => 69 , p => False), (a => 125, b => 133, p => False), (a => 11 , b => 19 , p => False), (a => 27 , b => 35 , p => False), (a => 43 , b => 51 , p => False), (a => 59 , b => 67 , p => False), (a => 75 , b => 83 , p => False), (a => 123, b => 131, p => False), (a => 139, b => 147, p => False), (a => 15 , b => 23 , p => False), (a => 31 , b => 39 , p => False), (a => 63 , b => 71 , p => False), (a => 127, b => 135, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 44 , b => 343, p => True ), (a => 45 , b => 342, p => True ), (a => 46 , b => 341, p => True ), (a => 47 , b => 340, p => True ), (a => 52 , b => 339, p => True ), (a => 53 , b => 338, p => True ), (a => 54 , b => 337, p => True ), (a => 55 , b => 336, p => True ), (a => 76 , b => 335, p => True ), (a => 77 , b => 334, p => True ), (a => 78 , b => 333, p => True ), (a => 79 , b => 332, p => True ), (a => 84 , b => 331, p => True ), (a => 85 , b => 330, p => True ), (a => 86 , b => 329, p => True ), (a => 87 , b => 328, p => True ), (a => 88 , b => 327, p => True ), (a => 89 , b => 326, p => True ), (a => 90 , b => 325, p => True ), (a => 91 , b => 324, p => True ), (a => 92 , b => 323, p => True ), (a => 93 , b => 322, p => True ), (a => 94 , b => 321, p => True ), (a => 95 , b => 320, p => True ), (a => 96 , b => 319, p => True ), (a => 97 , b => 318, p => True ), (a => 98 , b => 317, p => True ), (a => 99 , b => 316, p => True ), (a => 100, b => 315, p => True ), (a => 101, b => 314, p => True ), (a => 102, b => 313, p => True ), (a => 103, b => 312, p => True ), (a => 104, b => 311, p => True ), (a => 105, b => 310, p => True ), (a => 106, b => 309, p => True ), (a => 107, b => 308, p => True ), (a => 108, b => 307, p => True ), (a => 109, b => 306, p => True ), (a => 110, b => 305, p => True ), (a => 111, b => 304, p => True ), (a => 112, b => 303, p => True ), (a => 113, b => 302, p => True ), (a => 114, b => 301, p => True ), (a => 115, b => 300, p => True ), (a => 116, b => 299, p => True ), (a => 117, b => 298, p => True ), (a => 118, b => 297, p => True ), (a => 119, b => 296, p => True ), (a => 140, b => 295, p => True ), (a => 141, b => 294, p => True ), (a => 142, b => 293, p => True ), (a => 143, b => 292, p => True ), (a => 148, b => 291, p => True ), (a => 149, b => 290, p => True ), (a => 150, b => 289, p => True ), (a => 151, b => 288, p => True ), (a => 152, b => 287, p => True ), (a => 153, b => 286, p => True ), (a => 154, b => 285, p => True ), (a => 155, b => 284, p => True ), (a => 156, b => 283, p => True ), (a => 157, b => 282, p => True ), (a => 158, b => 281, p => True ), (a => 159, b => 280, p => True ), (a => 160, b => 279, p => True ), (a => 161, b => 278, p => True ), (a => 162, b => 277, p => True ), (a => 163, b => 276, p => True ), (a => 164, b => 275, p => True ), (a => 165, b => 274, p => True ), (a => 166, b => 273, p => True ), (a => 167, b => 272, p => True ), (a => 168, b => 271, p => True ), (a => 169, b => 270, p => True ), (a => 170, b => 269, p => True ), (a => 171, b => 268, p => True ), (a => 172, b => 267, p => True ), (a => 173, b => 266, p => True ), (a => 174, b => 265, p => True ), (a => 175, b => 264, p => True ), (a => 176, b => 263, p => True ), (a => 177, b => 262, p => True ), (a => 178, b => 261, p => True ), (a => 179, b => 260, p => True ), (a => 180, b => 259, p => True ), (a => 181, b => 258, p => True ), (a => 182, b => 257, p => True ), (a => 183, b => 256, p => True ), (a => 184, b => 255, p => True ), (a => 185, b => 254, p => True ), (a => 186, b => 253, p => True ), (a => 187, b => 252, p => True ), (a => 188, b => 251, p => True ), (a => 189, b => 250, p => True ), (a => 190, b => 249, p => True ), (a => 191, b => 248, p => True ), (a => 192, b => 247, p => True ), (a => 193, b => 246, p => True ), (a => 194, b => 245, p => True ), (a => 195, b => 244, p => True ), (a => 196, b => 243, p => True ), (a => 197, b => 242, p => True ), (a => 198, b => 241, p => True ), (a => 199, b => 240, p => True ), (a => 200, b => 239, p => True ), (a => 201, b => 238, p => True ), (a => 202, b => 237, p => True ), (a => 203, b => 236, p => True ), (a => 204, b => 235, p => True ), (a => 205, b => 234, p => True ), (a => 206, b => 233, p => True ), (a => 207, b => 232, p => True ), (a => 208, b => 231, p => True ), (a => 209, b => 230, p => True ), (a => 210, b => 229, p => True ), (a => 211, b => 228, p => True ), (a => 212, b => 227, p => True ), (a => 213, b => 226, p => True ), (a => 214, b => 225, p => True ), (a => 215, b => 224, p => True ), (a => 216, b => 223, p => True ), (a => 217, b => 222, p => True ), (a => 218, b => 221, p => True ), (a => 219, b => 220, p => True )),
                    ((a => 4  , b => 8  , p => False), (a => 12 , b => 16 , p => False), (a => 20 , b => 24 , p => False), (a => 28 , b => 32 , p => False), (a => 36 , b => 40 , p => False), (a => 60 , b => 64 , p => False), (a => 68 , b => 72 , p => False), (a => 124, b => 128, p => False), (a => 132, b => 136, p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 22 , b => 26 , p => False), (a => 30 , b => 34 , p => False), (a => 38 , b => 42 , p => False), (a => 62 , b => 66 , p => False), (a => 70 , b => 74 , p => False), (a => 126, b => 130, p => False), (a => 134, b => 138, p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 21 , b => 25 , p => False), (a => 29 , b => 33 , p => False), (a => 37 , b => 41 , p => False), (a => 61 , b => 65 , p => False), (a => 69 , b => 73 , p => False), (a => 125, b => 129, p => False), (a => 133, b => 137, p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 23 , b => 27 , p => False), (a => 31 , b => 35 , p => False), (a => 39 , b => 43 , p => False), (a => 63 , b => 67 , p => False), (a => 71 , b => 75 , p => False), (a => 127, b => 131, p => False), (a => 135, b => 139, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 44 , b => 347, p => True ), (a => 45 , b => 346, p => True ), (a => 46 , b => 345, p => True ), (a => 47 , b => 344, p => True ), (a => 48 , b => 343, p => True ), (a => 49 , b => 342, p => True ), (a => 50 , b => 341, p => True ), (a => 51 , b => 340, p => True ), (a => 52 , b => 339, p => True ), (a => 53 , b => 338, p => True ), (a => 54 , b => 337, p => True ), (a => 55 , b => 336, p => True ), (a => 56 , b => 335, p => True ), (a => 57 , b => 334, p => True ), (a => 58 , b => 333, p => True ), (a => 59 , b => 332, p => True ), (a => 76 , b => 331, p => True ), (a => 77 , b => 330, p => True ), (a => 78 , b => 329, p => True ), (a => 79 , b => 328, p => True ), (a => 80 , b => 327, p => True ), (a => 81 , b => 326, p => True ), (a => 82 , b => 325, p => True ), (a => 83 , b => 324, p => True ), (a => 84 , b => 323, p => True ), (a => 85 , b => 322, p => True ), (a => 86 , b => 321, p => True ), (a => 87 , b => 320, p => True ), (a => 88 , b => 319, p => True ), (a => 89 , b => 318, p => True ), (a => 90 , b => 317, p => True ), (a => 91 , b => 316, p => True ), (a => 92 , b => 315, p => True ), (a => 93 , b => 314, p => True ), (a => 94 , b => 313, p => True ), (a => 95 , b => 312, p => True ), (a => 96 , b => 311, p => True ), (a => 97 , b => 310, p => True ), (a => 98 , b => 309, p => True ), (a => 99 , b => 308, p => True ), (a => 100, b => 307, p => True ), (a => 101, b => 306, p => True ), (a => 102, b => 305, p => True ), (a => 103, b => 304, p => True ), (a => 104, b => 303, p => True ), (a => 105, b => 302, p => True ), (a => 106, b => 301, p => True ), (a => 107, b => 300, p => True ), (a => 108, b => 299, p => True ), (a => 109, b => 298, p => True ), (a => 110, b => 297, p => True ), (a => 111, b => 296, p => True ), (a => 112, b => 295, p => True ), (a => 113, b => 294, p => True ), (a => 114, b => 293, p => True ), (a => 115, b => 292, p => True ), (a => 116, b => 291, p => True ), (a => 117, b => 290, p => True ), (a => 118, b => 289, p => True ), (a => 119, b => 288, p => True ), (a => 120, b => 287, p => True ), (a => 121, b => 286, p => True ), (a => 122, b => 285, p => True ), (a => 123, b => 284, p => True ), (a => 140, b => 283, p => True ), (a => 141, b => 282, p => True ), (a => 142, b => 281, p => True ), (a => 143, b => 280, p => True ), (a => 144, b => 279, p => True ), (a => 145, b => 278, p => True ), (a => 146, b => 277, p => True ), (a => 147, b => 276, p => True ), (a => 148, b => 275, p => True ), (a => 149, b => 274, p => True ), (a => 150, b => 273, p => True ), (a => 151, b => 272, p => True ), (a => 152, b => 271, p => True ), (a => 153, b => 270, p => True ), (a => 154, b => 269, p => True ), (a => 155, b => 268, p => True ), (a => 156, b => 267, p => True ), (a => 157, b => 266, p => True ), (a => 158, b => 265, p => True ), (a => 159, b => 264, p => True ), (a => 160, b => 263, p => True ), (a => 161, b => 262, p => True ), (a => 162, b => 261, p => True ), (a => 163, b => 260, p => True ), (a => 164, b => 259, p => True ), (a => 165, b => 258, p => True ), (a => 166, b => 257, p => True ), (a => 167, b => 256, p => True ), (a => 168, b => 255, p => True ), (a => 169, b => 254, p => True ), (a => 170, b => 253, p => True ), (a => 171, b => 252, p => True ), (a => 172, b => 251, p => True ), (a => 173, b => 250, p => True ), (a => 174, b => 249, p => True ), (a => 175, b => 248, p => True ), (a => 176, b => 247, p => True ), (a => 177, b => 246, p => True ), (a => 178, b => 245, p => True ), (a => 179, b => 244, p => True ), (a => 180, b => 243, p => True ), (a => 181, b => 242, p => True ), (a => 182, b => 241, p => True ), (a => 183, b => 240, p => True ), (a => 184, b => 239, p => True ), (a => 185, b => 238, p => True ), (a => 186, b => 237, p => True ), (a => 187, b => 236, p => True ), (a => 188, b => 235, p => True ), (a => 189, b => 234, p => True ), (a => 190, b => 233, p => True ), (a => 191, b => 232, p => True ), (a => 192, b => 231, p => True ), (a => 193, b => 230, p => True ), (a => 194, b => 229, p => True ), (a => 195, b => 228, p => True ), (a => 196, b => 227, p => True ), (a => 197, b => 226, p => True ), (a => 198, b => 225, p => True ), (a => 199, b => 224, p => True ), (a => 200, b => 223, p => True ), (a => 201, b => 222, p => True ), (a => 202, b => 221, p => True ), (a => 203, b => 220, p => True ), (a => 204, b => 219, p => True ), (a => 205, b => 218, p => True ), (a => 206, b => 217, p => True ), (a => 207, b => 216, p => True ), (a => 208, b => 215, p => True ), (a => 209, b => 214, p => True ), (a => 210, b => 213, p => True ), (a => 211, b => 212, p => True )),
                    ((a => 2  , b => 4  , p => False), (a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 18 , b => 20 , p => False), (a => 22 , b => 24 , p => False), (a => 30 , b => 32 , p => False), (a => 34 , b => 36 , p => False), (a => 38 , b => 40 , p => False), (a => 62 , b => 64 , p => False), (a => 66 , b => 68 , p => False), (a => 70 , b => 72 , p => False), (a => 126, b => 128, p => False), (a => 130, b => 132, p => False), (a => 134, b => 136, p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 19 , b => 21 , p => False), (a => 23 , b => 25 , p => False), (a => 31 , b => 33 , p => False), (a => 35 , b => 37 , p => False), (a => 39 , b => 41 , p => False), (a => 63 , b => 65 , p => False), (a => 67 , b => 69 , p => False), (a => 71 , b => 73 , p => False), (a => 127, b => 129, p => False), (a => 131, b => 133, p => False), (a => 135, b => 137, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 26 , b => 349, p => True ), (a => 27 , b => 348, p => True ), (a => 28 , b => 347, p => True ), (a => 29 , b => 346, p => True ), (a => 42 , b => 345, p => True ), (a => 43 , b => 344, p => True ), (a => 44 , b => 343, p => True ), (a => 45 , b => 342, p => True ), (a => 46 , b => 341, p => True ), (a => 47 , b => 340, p => True ), (a => 48 , b => 339, p => True ), (a => 49 , b => 338, p => True ), (a => 50 , b => 337, p => True ), (a => 51 , b => 336, p => True ), (a => 52 , b => 335, p => True ), (a => 53 , b => 334, p => True ), (a => 54 , b => 333, p => True ), (a => 55 , b => 332, p => True ), (a => 56 , b => 331, p => True ), (a => 57 , b => 330, p => True ), (a => 58 , b => 329, p => True ), (a => 59 , b => 328, p => True ), (a => 60 , b => 327, p => True ), (a => 61 , b => 326, p => True ), (a => 74 , b => 325, p => True ), (a => 75 , b => 324, p => True ), (a => 76 , b => 323, p => True ), (a => 77 , b => 322, p => True ), (a => 78 , b => 321, p => True ), (a => 79 , b => 320, p => True ), (a => 80 , b => 319, p => True ), (a => 81 , b => 318, p => True ), (a => 82 , b => 317, p => True ), (a => 83 , b => 316, p => True ), (a => 84 , b => 315, p => True ), (a => 85 , b => 314, p => True ), (a => 86 , b => 313, p => True ), (a => 87 , b => 312, p => True ), (a => 88 , b => 311, p => True ), (a => 89 , b => 310, p => True ), (a => 90 , b => 309, p => True ), (a => 91 , b => 308, p => True ), (a => 92 , b => 307, p => True ), (a => 93 , b => 306, p => True ), (a => 94 , b => 305, p => True ), (a => 95 , b => 304, p => True ), (a => 96 , b => 303, p => True ), (a => 97 , b => 302, p => True ), (a => 98 , b => 301, p => True ), (a => 99 , b => 300, p => True ), (a => 100, b => 299, p => True ), (a => 101, b => 298, p => True ), (a => 102, b => 297, p => True ), (a => 103, b => 296, p => True ), (a => 104, b => 295, p => True ), (a => 105, b => 294, p => True ), (a => 106, b => 293, p => True ), (a => 107, b => 292, p => True ), (a => 108, b => 291, p => True ), (a => 109, b => 290, p => True ), (a => 110, b => 289, p => True ), (a => 111, b => 288, p => True ), (a => 112, b => 287, p => True ), (a => 113, b => 286, p => True ), (a => 114, b => 285, p => True ), (a => 115, b => 284, p => True ), (a => 116, b => 283, p => True ), (a => 117, b => 282, p => True ), (a => 118, b => 281, p => True ), (a => 119, b => 280, p => True ), (a => 120, b => 279, p => True ), (a => 121, b => 278, p => True ), (a => 122, b => 277, p => True ), (a => 123, b => 276, p => True ), (a => 124, b => 275, p => True ), (a => 125, b => 274, p => True ), (a => 138, b => 273, p => True ), (a => 139, b => 272, p => True ), (a => 140, b => 271, p => True ), (a => 141, b => 270, p => True ), (a => 142, b => 269, p => True ), (a => 143, b => 268, p => True ), (a => 144, b => 267, p => True ), (a => 145, b => 266, p => True ), (a => 146, b => 265, p => True ), (a => 147, b => 264, p => True ), (a => 148, b => 263, p => True ), (a => 149, b => 262, p => True ), (a => 150, b => 261, p => True ), (a => 151, b => 260, p => True ), (a => 152, b => 259, p => True ), (a => 153, b => 258, p => True ), (a => 154, b => 257, p => True ), (a => 155, b => 256, p => True ), (a => 156, b => 255, p => True ), (a => 157, b => 254, p => True ), (a => 158, b => 253, p => True ), (a => 159, b => 252, p => True ), (a => 160, b => 251, p => True ), (a => 161, b => 250, p => True ), (a => 162, b => 249, p => True ), (a => 163, b => 248, p => True ), (a => 164, b => 247, p => True ), (a => 165, b => 246, p => True ), (a => 166, b => 245, p => True ), (a => 167, b => 244, p => True ), (a => 168, b => 243, p => True ), (a => 169, b => 242, p => True ), (a => 170, b => 241, p => True ), (a => 171, b => 240, p => True ), (a => 172, b => 239, p => True ), (a => 173, b => 238, p => True ), (a => 174, b => 237, p => True ), (a => 175, b => 236, p => True ), (a => 176, b => 235, p => True ), (a => 177, b => 234, p => True ), (a => 178, b => 233, p => True ), (a => 179, b => 232, p => True ), (a => 180, b => 231, p => True ), (a => 181, b => 230, p => True ), (a => 182, b => 229, p => True ), (a => 183, b => 228, p => True ), (a => 184, b => 227, p => True ), (a => 185, b => 226, p => True ), (a => 186, b => 225, p => True ), (a => 187, b => 224, p => True ), (a => 188, b => 223, p => True ), (a => 189, b => 222, p => True ), (a => 190, b => 221, p => True ), (a => 191, b => 220, p => True ), (a => 192, b => 219, p => True ), (a => 193, b => 218, p => True ), (a => 194, b => 217, p => True ), (a => 195, b => 216, p => True ), (a => 196, b => 215, p => True ), (a => 197, b => 214, p => True ), (a => 198, b => 213, p => True ), (a => 199, b => 212, p => True ), (a => 200, b => 211, p => True ), (a => 201, b => 210, p => True ), (a => 202, b => 209, p => True ), (a => 203, b => 208, p => True ), (a => 204, b => 207, p => True ), (a => 205, b => 206, p => True )),
                    ((a => 1  , b => 2  , p => False), (a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 17 , b => 18 , p => False), (a => 19 , b => 20 , p => False), (a => 21 , b => 22 , p => False), (a => 23 , b => 24 , p => False), (a => 31 , b => 32 , p => False), (a => 33 , b => 34 , p => False), (a => 35 , b => 36 , p => False), (a => 37 , b => 38 , p => False), (a => 39 , b => 40 , p => False), (a => 63 , b => 64 , p => False), (a => 65 , b => 66 , p => False), (a => 67 , b => 68 , p => False), (a => 69 , b => 70 , p => False), (a => 71 , b => 72 , p => False), (a => 127, b => 128, p => False), (a => 129, b => 130, p => False), (a => 131, b => 132, p => False), (a => 133, b => 134, p => False), (a => 135, b => 136, p => False), (a => 0  , b => 351, p => True ), (a => 25 , b => 350, p => True ), (a => 26 , b => 349, p => True ), (a => 27 , b => 348, p => True ), (a => 28 , b => 347, p => True ), (a => 29 , b => 346, p => True ), (a => 30 , b => 345, p => True ), (a => 41 , b => 344, p => True ), (a => 42 , b => 343, p => True ), (a => 43 , b => 342, p => True ), (a => 44 , b => 341, p => True ), (a => 45 , b => 340, p => True ), (a => 46 , b => 339, p => True ), (a => 47 , b => 338, p => True ), (a => 48 , b => 337, p => True ), (a => 49 , b => 336, p => True ), (a => 50 , b => 335, p => True ), (a => 51 , b => 334, p => True ), (a => 52 , b => 333, p => True ), (a => 53 , b => 332, p => True ), (a => 54 , b => 331, p => True ), (a => 55 , b => 330, p => True ), (a => 56 , b => 329, p => True ), (a => 57 , b => 328, p => True ), (a => 58 , b => 327, p => True ), (a => 59 , b => 326, p => True ), (a => 60 , b => 325, p => True ), (a => 61 , b => 324, p => True ), (a => 62 , b => 323, p => True ), (a => 73 , b => 322, p => True ), (a => 74 , b => 321, p => True ), (a => 75 , b => 320, p => True ), (a => 76 , b => 319, p => True ), (a => 77 , b => 318, p => True ), (a => 78 , b => 317, p => True ), (a => 79 , b => 316, p => True ), (a => 80 , b => 315, p => True ), (a => 81 , b => 314, p => True ), (a => 82 , b => 313, p => True ), (a => 83 , b => 312, p => True ), (a => 84 , b => 311, p => True ), (a => 85 , b => 310, p => True ), (a => 86 , b => 309, p => True ), (a => 87 , b => 308, p => True ), (a => 88 , b => 307, p => True ), (a => 89 , b => 306, p => True ), (a => 90 , b => 305, p => True ), (a => 91 , b => 304, p => True ), (a => 92 , b => 303, p => True ), (a => 93 , b => 302, p => True ), (a => 94 , b => 301, p => True ), (a => 95 , b => 300, p => True ), (a => 96 , b => 299, p => True ), (a => 97 , b => 298, p => True ), (a => 98 , b => 297, p => True ), (a => 99 , b => 296, p => True ), (a => 100, b => 295, p => True ), (a => 101, b => 294, p => True ), (a => 102, b => 293, p => True ), (a => 103, b => 292, p => True ), (a => 104, b => 291, p => True ), (a => 105, b => 290, p => True ), (a => 106, b => 289, p => True ), (a => 107, b => 288, p => True ), (a => 108, b => 287, p => True ), (a => 109, b => 286, p => True ), (a => 110, b => 285, p => True ), (a => 111, b => 284, p => True ), (a => 112, b => 283, p => True ), (a => 113, b => 282, p => True ), (a => 114, b => 281, p => True ), (a => 115, b => 280, p => True ), (a => 116, b => 279, p => True ), (a => 117, b => 278, p => True ), (a => 118, b => 277, p => True ), (a => 119, b => 276, p => True ), (a => 120, b => 275, p => True ), (a => 121, b => 274, p => True ), (a => 122, b => 273, p => True ), (a => 123, b => 272, p => True ), (a => 124, b => 271, p => True ), (a => 125, b => 270, p => True ), (a => 126, b => 269, p => True ), (a => 137, b => 268, p => True ), (a => 138, b => 267, p => True ), (a => 139, b => 266, p => True ), (a => 140, b => 265, p => True ), (a => 141, b => 264, p => True ), (a => 142, b => 263, p => True ), (a => 143, b => 262, p => True ), (a => 144, b => 261, p => True ), (a => 145, b => 260, p => True ), (a => 146, b => 259, p => True ), (a => 147, b => 258, p => True ), (a => 148, b => 257, p => True ), (a => 149, b => 256, p => True ), (a => 150, b => 255, p => True ), (a => 151, b => 254, p => True ), (a => 152, b => 253, p => True ), (a => 153, b => 252, p => True ), (a => 154, b => 251, p => True ), (a => 155, b => 250, p => True ), (a => 156, b => 249, p => True ), (a => 157, b => 248, p => True ), (a => 158, b => 247, p => True ), (a => 159, b => 246, p => True ), (a => 160, b => 245, p => True ), (a => 161, b => 244, p => True ), (a => 162, b => 243, p => True ), (a => 163, b => 242, p => True ), (a => 164, b => 241, p => True ), (a => 165, b => 240, p => True ), (a => 166, b => 239, p => True ), (a => 167, b => 238, p => True ), (a => 168, b => 237, p => True ), (a => 169, b => 236, p => True ), (a => 170, b => 235, p => True ), (a => 171, b => 234, p => True ), (a => 172, b => 233, p => True ), (a => 173, b => 232, p => True ), (a => 174, b => 231, p => True ), (a => 175, b => 230, p => True ), (a => 176, b => 229, p => True ), (a => 177, b => 228, p => True ), (a => 178, b => 227, p => True ), (a => 179, b => 226, p => True ), (a => 180, b => 225, p => True ), (a => 181, b => 224, p => True ), (a => 182, b => 223, p => True ), (a => 183, b => 222, p => True ), (a => 184, b => 221, p => True ), (a => 185, b => 220, p => True ), (a => 186, b => 219, p => True ), (a => 187, b => 218, p => True ), (a => 188, b => 217, p => True ), (a => 189, b => 216, p => True ), (a => 190, b => 215, p => True ), (a => 191, b => 214, p => True ), (a => 192, b => 213, p => True ), (a => 193, b => 212, p => True ), (a => 194, b => 211, p => True ), (a => 195, b => 210, p => True ), (a => 196, b => 209, p => True ), (a => 197, b => 208, p => True ), (a => 198, b => 207, p => True ), (a => 199, b => 206, p => True ), (a => 200, b => 205, p => True ), (a => 201, b => 204, p => True ), (a => 202, b => 203, p => True )),
                    ((a => 64 , b => 320, p => False), (a => 32 , b => 288, p => False), (a => 16 , b => 272, p => False), (a => 8  , b => 264, p => False), (a => 4  , b => 260, p => False), (a => 68 , b => 324, p => False), (a => 36 , b => 292, p => False), (a => 20 , b => 276, p => False), (a => 12 , b => 268, p => False), (a => 2  , b => 258, p => False), (a => 66 , b => 322, p => False), (a => 34 , b => 290, p => False), (a => 18 , b => 274, p => False), (a => 10 , b => 266, p => False), (a => 6  , b => 262, p => False), (a => 70 , b => 326, p => False), (a => 38 , b => 294, p => False), (a => 22 , b => 278, p => False), (a => 14 , b => 270, p => False), (a => 1  , b => 257, p => False), (a => 65 , b => 321, p => False), (a => 33 , b => 289, p => False), (a => 17 , b => 273, p => False), (a => 9  , b => 265, p => False), (a => 5  , b => 261, p => False), (a => 69 , b => 325, p => False), (a => 37 , b => 293, p => False), (a => 21 , b => 277, p => False), (a => 13 , b => 269, p => False), (a => 3  , b => 259, p => False), (a => 67 , b => 323, p => False), (a => 35 , b => 291, p => False), (a => 19 , b => 275, p => False), (a => 11 , b => 267, p => False), (a => 7  , b => 263, p => False), (a => 71 , b => 327, p => False), (a => 39 , b => 295, p => False), (a => 23 , b => 279, p => False), (a => 15 , b => 271, p => False), (a => 128, b => 256, p => False), (a => 0  , b => 351, p => True ), (a => 24 , b => 350, p => True ), (a => 25 , b => 349, p => True ), (a => 26 , b => 348, p => True ), (a => 27 , b => 347, p => True ), (a => 28 , b => 346, p => True ), (a => 29 , b => 345, p => True ), (a => 30 , b => 344, p => True ), (a => 31 , b => 343, p => True ), (a => 40 , b => 342, p => True ), (a => 41 , b => 341, p => True ), (a => 42 , b => 340, p => True ), (a => 43 , b => 339, p => True ), (a => 44 , b => 338, p => True ), (a => 45 , b => 337, p => True ), (a => 46 , b => 336, p => True ), (a => 47 , b => 335, p => True ), (a => 48 , b => 334, p => True ), (a => 49 , b => 333, p => True ), (a => 50 , b => 332, p => True ), (a => 51 , b => 331, p => True ), (a => 52 , b => 330, p => True ), (a => 53 , b => 329, p => True ), (a => 54 , b => 328, p => True ), (a => 55 , b => 319, p => True ), (a => 56 , b => 318, p => True ), (a => 57 , b => 317, p => True ), (a => 58 , b => 316, p => True ), (a => 59 , b => 315, p => True ), (a => 60 , b => 314, p => True ), (a => 61 , b => 313, p => True ), (a => 62 , b => 312, p => True ), (a => 63 , b => 311, p => True ), (a => 72 , b => 310, p => True ), (a => 73 , b => 309, p => True ), (a => 74 , b => 308, p => True ), (a => 75 , b => 307, p => True ), (a => 76 , b => 306, p => True ), (a => 77 , b => 305, p => True ), (a => 78 , b => 304, p => True ), (a => 79 , b => 303, p => True ), (a => 80 , b => 302, p => True ), (a => 81 , b => 301, p => True ), (a => 82 , b => 300, p => True ), (a => 83 , b => 299, p => True ), (a => 84 , b => 298, p => True ), (a => 85 , b => 297, p => True ), (a => 86 , b => 296, p => True ), (a => 87 , b => 287, p => True ), (a => 88 , b => 286, p => True ), (a => 89 , b => 285, p => True ), (a => 90 , b => 284, p => True ), (a => 91 , b => 283, p => True ), (a => 92 , b => 282, p => True ), (a => 93 , b => 281, p => True ), (a => 94 , b => 280, p => True ), (a => 95 , b => 255, p => True ), (a => 96 , b => 254, p => True ), (a => 97 , b => 253, p => True ), (a => 98 , b => 252, p => True ), (a => 99 , b => 251, p => True ), (a => 100, b => 250, p => True ), (a => 101, b => 249, p => True ), (a => 102, b => 248, p => True ), (a => 103, b => 247, p => True ), (a => 104, b => 246, p => True ), (a => 105, b => 245, p => True ), (a => 106, b => 244, p => True ), (a => 107, b => 243, p => True ), (a => 108, b => 242, p => True ), (a => 109, b => 241, p => True ), (a => 110, b => 240, p => True ), (a => 111, b => 239, p => True ), (a => 112, b => 238, p => True ), (a => 113, b => 237, p => True ), (a => 114, b => 236, p => True ), (a => 115, b => 235, p => True ), (a => 116, b => 234, p => True ), (a => 117, b => 233, p => True ), (a => 118, b => 232, p => True ), (a => 119, b => 231, p => True ), (a => 120, b => 230, p => True ), (a => 121, b => 229, p => True ), (a => 122, b => 228, p => True ), (a => 123, b => 227, p => True ), (a => 124, b => 226, p => True ), (a => 125, b => 225, p => True ), (a => 126, b => 224, p => True ), (a => 127, b => 223, p => True ), (a => 129, b => 222, p => True ), (a => 130, b => 221, p => True ), (a => 131, b => 220, p => True ), (a => 132, b => 219, p => True ), (a => 133, b => 218, p => True ), (a => 134, b => 217, p => True ), (a => 135, b => 216, p => True ), (a => 136, b => 215, p => True ), (a => 137, b => 214, p => True ), (a => 138, b => 213, p => True ), (a => 139, b => 212, p => True ), (a => 140, b => 211, p => True ), (a => 141, b => 210, p => True ), (a => 142, b => 209, p => True ), (a => 143, b => 208, p => True ), (a => 144, b => 207, p => True ), (a => 145, b => 206, p => True ), (a => 146, b => 205, p => True ), (a => 147, b => 204, p => True ), (a => 148, b => 203, p => True ), (a => 149, b => 202, p => True ), (a => 150, b => 201, p => True ), (a => 151, b => 200, p => True ), (a => 152, b => 199, p => True ), (a => 153, b => 198, p => True ), (a => 154, b => 197, p => True ), (a => 155, b => 196, p => True ), (a => 156, b => 195, p => True ), (a => 157, b => 194, p => True ), (a => 158, b => 193, p => True ), (a => 159, b => 192, p => True ), (a => 160, b => 191, p => True ), (a => 161, b => 190, p => True ), (a => 162, b => 189, p => True ), (a => 163, b => 188, p => True ), (a => 164, b => 187, p => True ), (a => 165, b => 186, p => True ), (a => 166, b => 185, p => True ), (a => 167, b => 184, p => True ), (a => 168, b => 183, p => True ), (a => 169, b => 182, p => True ), (a => 170, b => 181, p => True ), (a => 171, b => 180, p => True ), (a => 172, b => 179, p => True ), (a => 173, b => 178, p => True ), (a => 174, b => 177, p => True ), (a => 175, b => 176, p => True )),
                    ((a => 132, b => 260, p => False), (a => 130, b => 258, p => False), (a => 134, b => 262, p => False), (a => 129, b => 257, p => False), (a => 133, b => 261, p => False), (a => 131, b => 259, p => False), (a => 135, b => 263, p => False), (a => 64 , b => 128, p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 343, p => True ), (a => 9  , b => 342, p => True ), (a => 10 , b => 341, p => True ), (a => 11 , b => 340, p => True ), (a => 12 , b => 339, p => True ), (a => 13 , b => 338, p => True ), (a => 14 , b => 337, p => True ), (a => 15 , b => 336, p => True ), (a => 16 , b => 335, p => True ), (a => 17 , b => 334, p => True ), (a => 18 , b => 333, p => True ), (a => 19 , b => 332, p => True ), (a => 20 , b => 331, p => True ), (a => 21 , b => 330, p => True ), (a => 22 , b => 329, p => True ), (a => 23 , b => 328, p => True ), (a => 24 , b => 327, p => True ), (a => 25 , b => 326, p => True ), (a => 26 , b => 325, p => True ), (a => 27 , b => 324, p => True ), (a => 28 , b => 323, p => True ), (a => 29 , b => 322, p => True ), (a => 30 , b => 321, p => True ), (a => 31 , b => 320, p => True ), (a => 32 , b => 319, p => True ), (a => 33 , b => 318, p => True ), (a => 34 , b => 317, p => True ), (a => 35 , b => 316, p => True ), (a => 36 , b => 315, p => True ), (a => 37 , b => 314, p => True ), (a => 38 , b => 313, p => True ), (a => 39 , b => 312, p => True ), (a => 40 , b => 311, p => True ), (a => 41 , b => 310, p => True ), (a => 42 , b => 309, p => True ), (a => 43 , b => 308, p => True ), (a => 44 , b => 307, p => True ), (a => 45 , b => 306, p => True ), (a => 46 , b => 305, p => True ), (a => 47 , b => 304, p => True ), (a => 48 , b => 303, p => True ), (a => 49 , b => 302, p => True ), (a => 50 , b => 301, p => True ), (a => 51 , b => 300, p => True ), (a => 52 , b => 299, p => True ), (a => 53 , b => 298, p => True ), (a => 54 , b => 297, p => True ), (a => 55 , b => 296, p => True ), (a => 56 , b => 295, p => True ), (a => 57 , b => 294, p => True ), (a => 58 , b => 293, p => True ), (a => 59 , b => 292, p => True ), (a => 60 , b => 291, p => True ), (a => 61 , b => 290, p => True ), (a => 62 , b => 289, p => True ), (a => 63 , b => 288, p => True ), (a => 65 , b => 287, p => True ), (a => 66 , b => 286, p => True ), (a => 67 , b => 285, p => True ), (a => 68 , b => 284, p => True ), (a => 69 , b => 283, p => True ), (a => 70 , b => 282, p => True ), (a => 71 , b => 281, p => True ), (a => 72 , b => 280, p => True ), (a => 73 , b => 279, p => True ), (a => 74 , b => 278, p => True ), (a => 75 , b => 277, p => True ), (a => 76 , b => 276, p => True ), (a => 77 , b => 275, p => True ), (a => 78 , b => 274, p => True ), (a => 79 , b => 273, p => True ), (a => 80 , b => 272, p => True ), (a => 81 , b => 271, p => True ), (a => 82 , b => 270, p => True ), (a => 83 , b => 269, p => True ), (a => 84 , b => 268, p => True ), (a => 85 , b => 267, p => True ), (a => 86 , b => 266, p => True ), (a => 87 , b => 265, p => True ), (a => 88 , b => 264, p => True ), (a => 89 , b => 256, p => True ), (a => 90 , b => 255, p => True ), (a => 91 , b => 254, p => True ), (a => 92 , b => 253, p => True ), (a => 93 , b => 252, p => True ), (a => 94 , b => 251, p => True ), (a => 95 , b => 250, p => True ), (a => 96 , b => 249, p => True ), (a => 97 , b => 248, p => True ), (a => 98 , b => 247, p => True ), (a => 99 , b => 246, p => True ), (a => 100, b => 245, p => True ), (a => 101, b => 244, p => True ), (a => 102, b => 243, p => True ), (a => 103, b => 242, p => True ), (a => 104, b => 241, p => True ), (a => 105, b => 240, p => True ), (a => 106, b => 239, p => True ), (a => 107, b => 238, p => True ), (a => 108, b => 237, p => True ), (a => 109, b => 236, p => True ), (a => 110, b => 235, p => True ), (a => 111, b => 234, p => True ), (a => 112, b => 233, p => True ), (a => 113, b => 232, p => True ), (a => 114, b => 231, p => True ), (a => 115, b => 230, p => True ), (a => 116, b => 229, p => True ), (a => 117, b => 228, p => True ), (a => 118, b => 227, p => True ), (a => 119, b => 226, p => True ), (a => 120, b => 225, p => True ), (a => 121, b => 224, p => True ), (a => 122, b => 223, p => True ), (a => 123, b => 222, p => True ), (a => 124, b => 221, p => True ), (a => 125, b => 220, p => True ), (a => 126, b => 219, p => True ), (a => 127, b => 218, p => True ), (a => 136, b => 217, p => True ), (a => 137, b => 216, p => True ), (a => 138, b => 215, p => True ), (a => 139, b => 214, p => True ), (a => 140, b => 213, p => True ), (a => 141, b => 212, p => True ), (a => 142, b => 211, p => True ), (a => 143, b => 210, p => True ), (a => 144, b => 209, p => True ), (a => 145, b => 208, p => True ), (a => 146, b => 207, p => True ), (a => 147, b => 206, p => True ), (a => 148, b => 205, p => True ), (a => 149, b => 204, p => True ), (a => 150, b => 203, p => True ), (a => 151, b => 202, p => True ), (a => 152, b => 201, p => True ), (a => 153, b => 200, p => True ), (a => 154, b => 199, p => True ), (a => 155, b => 198, p => True ), (a => 156, b => 197, p => True ), (a => 157, b => 196, p => True ), (a => 158, b => 195, p => True ), (a => 159, b => 194, p => True ), (a => 160, b => 193, p => True ), (a => 161, b => 192, p => True ), (a => 162, b => 191, p => True ), (a => 163, b => 190, p => True ), (a => 164, b => 189, p => True ), (a => 165, b => 188, p => True ), (a => 166, b => 187, p => True ), (a => 167, b => 186, p => True ), (a => 168, b => 185, p => True ), (a => 169, b => 184, p => True ), (a => 170, b => 183, p => True ), (a => 171, b => 182, p => True ), (a => 172, b => 181, p => True ), (a => 173, b => 180, p => True ), (a => 174, b => 179, p => True ), (a => 175, b => 178, p => True ), (a => 176, b => 177, p => True )),
                    ((a => 68 , b => 132, p => False), (a => 66 , b => 130, p => False), (a => 70 , b => 134, p => False), (a => 65 , b => 129, p => False), (a => 69 , b => 133, p => False), (a => 67 , b => 131, p => False), (a => 71 , b => 135, p => False), (a => 32 , b => 64 , p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 343, p => True ), (a => 9  , b => 342, p => True ), (a => 10 , b => 341, p => True ), (a => 11 , b => 340, p => True ), (a => 12 , b => 339, p => True ), (a => 13 , b => 338, p => True ), (a => 14 , b => 337, p => True ), (a => 15 , b => 336, p => True ), (a => 16 , b => 335, p => True ), (a => 17 , b => 334, p => True ), (a => 18 , b => 333, p => True ), (a => 19 , b => 332, p => True ), (a => 20 , b => 331, p => True ), (a => 21 , b => 330, p => True ), (a => 22 , b => 329, p => True ), (a => 23 , b => 328, p => True ), (a => 24 , b => 327, p => True ), (a => 25 , b => 326, p => True ), (a => 26 , b => 325, p => True ), (a => 27 , b => 324, p => True ), (a => 28 , b => 323, p => True ), (a => 29 , b => 322, p => True ), (a => 30 , b => 321, p => True ), (a => 31 , b => 320, p => True ), (a => 33 , b => 319, p => True ), (a => 34 , b => 318, p => True ), (a => 35 , b => 317, p => True ), (a => 36 , b => 316, p => True ), (a => 37 , b => 315, p => True ), (a => 38 , b => 314, p => True ), (a => 39 , b => 313, p => True ), (a => 40 , b => 312, p => True ), (a => 41 , b => 311, p => True ), (a => 42 , b => 310, p => True ), (a => 43 , b => 309, p => True ), (a => 44 , b => 308, p => True ), (a => 45 , b => 307, p => True ), (a => 46 , b => 306, p => True ), (a => 47 , b => 305, p => True ), (a => 48 , b => 304, p => True ), (a => 49 , b => 303, p => True ), (a => 50 , b => 302, p => True ), (a => 51 , b => 301, p => True ), (a => 52 , b => 300, p => True ), (a => 53 , b => 299, p => True ), (a => 54 , b => 298, p => True ), (a => 55 , b => 297, p => True ), (a => 56 , b => 296, p => True ), (a => 57 , b => 295, p => True ), (a => 58 , b => 294, p => True ), (a => 59 , b => 293, p => True ), (a => 60 , b => 292, p => True ), (a => 61 , b => 291, p => True ), (a => 62 , b => 290, p => True ), (a => 63 , b => 289, p => True ), (a => 72 , b => 288, p => True ), (a => 73 , b => 287, p => True ), (a => 74 , b => 286, p => True ), (a => 75 , b => 285, p => True ), (a => 76 , b => 284, p => True ), (a => 77 , b => 283, p => True ), (a => 78 , b => 282, p => True ), (a => 79 , b => 281, p => True ), (a => 80 , b => 280, p => True ), (a => 81 , b => 279, p => True ), (a => 82 , b => 278, p => True ), (a => 83 , b => 277, p => True ), (a => 84 , b => 276, p => True ), (a => 85 , b => 275, p => True ), (a => 86 , b => 274, p => True ), (a => 87 , b => 273, p => True ), (a => 88 , b => 272, p => True ), (a => 89 , b => 271, p => True ), (a => 90 , b => 270, p => True ), (a => 91 , b => 269, p => True ), (a => 92 , b => 268, p => True ), (a => 93 , b => 267, p => True ), (a => 94 , b => 266, p => True ), (a => 95 , b => 265, p => True ), (a => 96 , b => 264, p => True ), (a => 97 , b => 263, p => True ), (a => 98 , b => 262, p => True ), (a => 99 , b => 261, p => True ), (a => 100, b => 260, p => True ), (a => 101, b => 259, p => True ), (a => 102, b => 258, p => True ), (a => 103, b => 257, p => True ), (a => 104, b => 256, p => True ), (a => 105, b => 255, p => True ), (a => 106, b => 254, p => True ), (a => 107, b => 253, p => True ), (a => 108, b => 252, p => True ), (a => 109, b => 251, p => True ), (a => 110, b => 250, p => True ), (a => 111, b => 249, p => True ), (a => 112, b => 248, p => True ), (a => 113, b => 247, p => True ), (a => 114, b => 246, p => True ), (a => 115, b => 245, p => True ), (a => 116, b => 244, p => True ), (a => 117, b => 243, p => True ), (a => 118, b => 242, p => True ), (a => 119, b => 241, p => True ), (a => 120, b => 240, p => True ), (a => 121, b => 239, p => True ), (a => 122, b => 238, p => True ), (a => 123, b => 237, p => True ), (a => 124, b => 236, p => True ), (a => 125, b => 235, p => True ), (a => 126, b => 234, p => True ), (a => 127, b => 233, p => True ), (a => 128, b => 232, p => True ), (a => 136, b => 231, p => True ), (a => 137, b => 230, p => True ), (a => 138, b => 229, p => True ), (a => 139, b => 228, p => True ), (a => 140, b => 227, p => True ), (a => 141, b => 226, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 146, b => 221, p => True ), (a => 147, b => 220, p => True ), (a => 148, b => 219, p => True ), (a => 149, b => 218, p => True ), (a => 150, b => 217, p => True ), (a => 151, b => 216, p => True ), (a => 152, b => 215, p => True ), (a => 153, b => 214, p => True ), (a => 154, b => 213, p => True ), (a => 155, b => 212, p => True ), (a => 156, b => 211, p => True ), (a => 157, b => 210, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 162, b => 205, p => True ), (a => 163, b => 204, p => True ), (a => 164, b => 203, p => True ), (a => 165, b => 202, p => True ), (a => 166, b => 201, p => True ), (a => 167, b => 200, p => True ), (a => 168, b => 199, p => True ), (a => 169, b => 198, p => True ), (a => 170, b => 197, p => True ), (a => 171, b => 196, p => True ), (a => 172, b => 195, p => True ), (a => 173, b => 194, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True ), (a => 178, b => 189, p => True ), (a => 179, b => 188, p => True ), (a => 180, b => 187, p => True ), (a => 181, b => 186, p => True ), (a => 182, b => 185, p => True ), (a => 183, b => 184, p => True )),
                    ((a => 36 , b => 68 , p => False), (a => 34 , b => 66 , p => False), (a => 38 , b => 70 , p => False), (a => 33 , b => 65 , p => False), (a => 37 , b => 69 , p => False), (a => 35 , b => 67 , p => False), (a => 39 , b => 71 , p => False), (a => 16 , b => 32 , p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 8  , b => 343, p => True ), (a => 9  , b => 342, p => True ), (a => 10 , b => 341, p => True ), (a => 11 , b => 340, p => True ), (a => 12 , b => 339, p => True ), (a => 13 , b => 338, p => True ), (a => 14 , b => 337, p => True ), (a => 15 , b => 336, p => True ), (a => 17 , b => 335, p => True ), (a => 18 , b => 334, p => True ), (a => 19 , b => 333, p => True ), (a => 20 , b => 332, p => True ), (a => 21 , b => 331, p => True ), (a => 22 , b => 330, p => True ), (a => 23 , b => 329, p => True ), (a => 24 , b => 328, p => True ), (a => 25 , b => 327, p => True ), (a => 26 , b => 326, p => True ), (a => 27 , b => 325, p => True ), (a => 28 , b => 324, p => True ), (a => 29 , b => 323, p => True ), (a => 30 , b => 322, p => True ), (a => 31 , b => 321, p => True ), (a => 40 , b => 320, p => True ), (a => 41 , b => 319, p => True ), (a => 42 , b => 318, p => True ), (a => 43 , b => 317, p => True ), (a => 44 , b => 316, p => True ), (a => 45 , b => 315, p => True ), (a => 46 , b => 314, p => True ), (a => 47 , b => 313, p => True ), (a => 48 , b => 312, p => True ), (a => 49 , b => 311, p => True ), (a => 50 , b => 310, p => True ), (a => 51 , b => 309, p => True ), (a => 52 , b => 308, p => True ), (a => 53 , b => 307, p => True ), (a => 54 , b => 306, p => True ), (a => 55 , b => 305, p => True ), (a => 56 , b => 304, p => True ), (a => 57 , b => 303, p => True ), (a => 58 , b => 302, p => True ), (a => 59 , b => 301, p => True ), (a => 60 , b => 300, p => True ), (a => 61 , b => 299, p => True ), (a => 62 , b => 298, p => True ), (a => 63 , b => 297, p => True ), (a => 64 , b => 296, p => True ), (a => 72 , b => 295, p => True ), (a => 73 , b => 294, p => True ), (a => 74 , b => 293, p => True ), (a => 75 , b => 292, p => True ), (a => 76 , b => 291, p => True ), (a => 77 , b => 290, p => True ), (a => 78 , b => 289, p => True ), (a => 79 , b => 288, p => True ), (a => 80 , b => 287, p => True ), (a => 81 , b => 286, p => True ), (a => 82 , b => 285, p => True ), (a => 83 , b => 284, p => True ), (a => 84 , b => 283, p => True ), (a => 85 , b => 282, p => True ), (a => 86 , b => 281, p => True ), (a => 87 , b => 280, p => True ), (a => 88 , b => 279, p => True ), (a => 89 , b => 278, p => True ), (a => 90 , b => 277, p => True ), (a => 91 , b => 276, p => True ), (a => 92 , b => 275, p => True ), (a => 93 , b => 274, p => True ), (a => 94 , b => 273, p => True ), (a => 95 , b => 272, p => True ), (a => 96 , b => 271, p => True ), (a => 97 , b => 270, p => True ), (a => 98 , b => 269, p => True ), (a => 99 , b => 268, p => True ), (a => 100, b => 267, p => True ), (a => 101, b => 266, p => True ), (a => 102, b => 265, p => True ), (a => 103, b => 264, p => True ), (a => 104, b => 263, p => True ), (a => 105, b => 262, p => True ), (a => 106, b => 261, p => True ), (a => 107, b => 260, p => True ), (a => 108, b => 259, p => True ), (a => 109, b => 258, p => True ), (a => 110, b => 257, p => True ), (a => 111, b => 256, p => True ), (a => 112, b => 255, p => True ), (a => 113, b => 254, p => True ), (a => 114, b => 253, p => True ), (a => 115, b => 252, p => True ), (a => 116, b => 251, p => True ), (a => 117, b => 250, p => True ), (a => 118, b => 249, p => True ), (a => 119, b => 248, p => True ), (a => 120, b => 247, p => True ), (a => 121, b => 246, p => True ), (a => 122, b => 245, p => True ), (a => 123, b => 244, p => True ), (a => 124, b => 243, p => True ), (a => 125, b => 242, p => True ), (a => 126, b => 241, p => True ), (a => 127, b => 240, p => True ), (a => 128, b => 239, p => True ), (a => 129, b => 238, p => True ), (a => 130, b => 237, p => True ), (a => 131, b => 236, p => True ), (a => 132, b => 235, p => True ), (a => 133, b => 234, p => True ), (a => 134, b => 233, p => True ), (a => 135, b => 232, p => True ), (a => 136, b => 231, p => True ), (a => 137, b => 230, p => True ), (a => 138, b => 229, p => True ), (a => 139, b => 228, p => True ), (a => 140, b => 227, p => True ), (a => 141, b => 226, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 146, b => 221, p => True ), (a => 147, b => 220, p => True ), (a => 148, b => 219, p => True ), (a => 149, b => 218, p => True ), (a => 150, b => 217, p => True ), (a => 151, b => 216, p => True ), (a => 152, b => 215, p => True ), (a => 153, b => 214, p => True ), (a => 154, b => 213, p => True ), (a => 155, b => 212, p => True ), (a => 156, b => 211, p => True ), (a => 157, b => 210, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 162, b => 205, p => True ), (a => 163, b => 204, p => True ), (a => 164, b => 203, p => True ), (a => 165, b => 202, p => True ), (a => 166, b => 201, p => True ), (a => 167, b => 200, p => True ), (a => 168, b => 199, p => True ), (a => 169, b => 198, p => True ), (a => 170, b => 197, p => True ), (a => 171, b => 196, p => True ), (a => 172, b => 195, p => True ), (a => 173, b => 194, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True ), (a => 178, b => 189, p => True ), (a => 179, b => 188, p => True ), (a => 180, b => 187, p => True ), (a => 181, b => 186, p => True ), (a => 182, b => 185, p => True ), (a => 183, b => 184, p => True )),
                    ((a => 20 , b => 36 , p => False), (a => 18 , b => 34 , p => False), (a => 22 , b => 38 , p => False), (a => 17 , b => 33 , p => False), (a => 21 , b => 37 , p => False), (a => 19 , b => 35 , p => False), (a => 23 , b => 39 , p => False), (a => 8  , b => 16 , p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 4  , b => 347, p => True ), (a => 5  , b => 346, p => True ), (a => 6  , b => 345, p => True ), (a => 7  , b => 344, p => True ), (a => 9  , b => 343, p => True ), (a => 10 , b => 342, p => True ), (a => 11 , b => 341, p => True ), (a => 12 , b => 340, p => True ), (a => 13 , b => 339, p => True ), (a => 14 , b => 338, p => True ), (a => 15 , b => 337, p => True ), (a => 24 , b => 336, p => True ), (a => 25 , b => 335, p => True ), (a => 26 , b => 334, p => True ), (a => 27 , b => 333, p => True ), (a => 28 , b => 332, p => True ), (a => 29 , b => 331, p => True ), (a => 30 , b => 330, p => True ), (a => 31 , b => 329, p => True ), (a => 32 , b => 328, p => True ), (a => 40 , b => 327, p => True ), (a => 41 , b => 326, p => True ), (a => 42 , b => 325, p => True ), (a => 43 , b => 324, p => True ), (a => 44 , b => 323, p => True ), (a => 45 , b => 322, p => True ), (a => 46 , b => 321, p => True ), (a => 47 , b => 320, p => True ), (a => 48 , b => 319, p => True ), (a => 49 , b => 318, p => True ), (a => 50 , b => 317, p => True ), (a => 51 , b => 316, p => True ), (a => 52 , b => 315, p => True ), (a => 53 , b => 314, p => True ), (a => 54 , b => 313, p => True ), (a => 55 , b => 312, p => True ), (a => 56 , b => 311, p => True ), (a => 57 , b => 310, p => True ), (a => 58 , b => 309, p => True ), (a => 59 , b => 308, p => True ), (a => 60 , b => 307, p => True ), (a => 61 , b => 306, p => True ), (a => 62 , b => 305, p => True ), (a => 63 , b => 304, p => True ), (a => 64 , b => 303, p => True ), (a => 65 , b => 302, p => True ), (a => 66 , b => 301, p => True ), (a => 67 , b => 300, p => True ), (a => 68 , b => 299, p => True ), (a => 69 , b => 298, p => True ), (a => 70 , b => 297, p => True ), (a => 71 , b => 296, p => True ), (a => 72 , b => 295, p => True ), (a => 73 , b => 294, p => True ), (a => 74 , b => 293, p => True ), (a => 75 , b => 292, p => True ), (a => 76 , b => 291, p => True ), (a => 77 , b => 290, p => True ), (a => 78 , b => 289, p => True ), (a => 79 , b => 288, p => True ), (a => 80 , b => 287, p => True ), (a => 81 , b => 286, p => True ), (a => 82 , b => 285, p => True ), (a => 83 , b => 284, p => True ), (a => 84 , b => 283, p => True ), (a => 85 , b => 282, p => True ), (a => 86 , b => 281, p => True ), (a => 87 , b => 280, p => True ), (a => 88 , b => 279, p => True ), (a => 89 , b => 278, p => True ), (a => 90 , b => 277, p => True ), (a => 91 , b => 276, p => True ), (a => 92 , b => 275, p => True ), (a => 93 , b => 274, p => True ), (a => 94 , b => 273, p => True ), (a => 95 , b => 272, p => True ), (a => 96 , b => 271, p => True ), (a => 97 , b => 270, p => True ), (a => 98 , b => 269, p => True ), (a => 99 , b => 268, p => True ), (a => 100, b => 267, p => True ), (a => 101, b => 266, p => True ), (a => 102, b => 265, p => True ), (a => 103, b => 264, p => True ), (a => 104, b => 263, p => True ), (a => 105, b => 262, p => True ), (a => 106, b => 261, p => True ), (a => 107, b => 260, p => True ), (a => 108, b => 259, p => True ), (a => 109, b => 258, p => True ), (a => 110, b => 257, p => True ), (a => 111, b => 256, p => True ), (a => 112, b => 255, p => True ), (a => 113, b => 254, p => True ), (a => 114, b => 253, p => True ), (a => 115, b => 252, p => True ), (a => 116, b => 251, p => True ), (a => 117, b => 250, p => True ), (a => 118, b => 249, p => True ), (a => 119, b => 248, p => True ), (a => 120, b => 247, p => True ), (a => 121, b => 246, p => True ), (a => 122, b => 245, p => True ), (a => 123, b => 244, p => True ), (a => 124, b => 243, p => True ), (a => 125, b => 242, p => True ), (a => 126, b => 241, p => True ), (a => 127, b => 240, p => True ), (a => 128, b => 239, p => True ), (a => 129, b => 238, p => True ), (a => 130, b => 237, p => True ), (a => 131, b => 236, p => True ), (a => 132, b => 235, p => True ), (a => 133, b => 234, p => True ), (a => 134, b => 233, p => True ), (a => 135, b => 232, p => True ), (a => 136, b => 231, p => True ), (a => 137, b => 230, p => True ), (a => 138, b => 229, p => True ), (a => 139, b => 228, p => True ), (a => 140, b => 227, p => True ), (a => 141, b => 226, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 146, b => 221, p => True ), (a => 147, b => 220, p => True ), (a => 148, b => 219, p => True ), (a => 149, b => 218, p => True ), (a => 150, b => 217, p => True ), (a => 151, b => 216, p => True ), (a => 152, b => 215, p => True ), (a => 153, b => 214, p => True ), (a => 154, b => 213, p => True ), (a => 155, b => 212, p => True ), (a => 156, b => 211, p => True ), (a => 157, b => 210, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 162, b => 205, p => True ), (a => 163, b => 204, p => True ), (a => 164, b => 203, p => True ), (a => 165, b => 202, p => True ), (a => 166, b => 201, p => True ), (a => 167, b => 200, p => True ), (a => 168, b => 199, p => True ), (a => 169, b => 198, p => True ), (a => 170, b => 197, p => True ), (a => 171, b => 196, p => True ), (a => 172, b => 195, p => True ), (a => 173, b => 194, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True ), (a => 178, b => 189, p => True ), (a => 179, b => 188, p => True ), (a => 180, b => 187, p => True ), (a => 181, b => 186, p => True ), (a => 182, b => 185, p => True ), (a => 183, b => 184, p => True )),
                    ((a => 12 , b => 20 , p => False), (a => 10 , b => 18 , p => False), (a => 14 , b => 22 , p => False), (a => 9  , b => 17 , p => False), (a => 13 , b => 21 , p => False), (a => 11 , b => 19 , p => False), (a => 15 , b => 23 , p => False), (a => 4  , b => 8  , p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 3  , b => 348, p => True ), (a => 5  , b => 347, p => True ), (a => 6  , b => 346, p => True ), (a => 7  , b => 345, p => True ), (a => 16 , b => 344, p => True ), (a => 24 , b => 343, p => True ), (a => 25 , b => 342, p => True ), (a => 26 , b => 341, p => True ), (a => 27 , b => 340, p => True ), (a => 28 , b => 339, p => True ), (a => 29 , b => 338, p => True ), (a => 30 , b => 337, p => True ), (a => 31 , b => 336, p => True ), (a => 32 , b => 335, p => True ), (a => 33 , b => 334, p => True ), (a => 34 , b => 333, p => True ), (a => 35 , b => 332, p => True ), (a => 36 , b => 331, p => True ), (a => 37 , b => 330, p => True ), (a => 38 , b => 329, p => True ), (a => 39 , b => 328, p => True ), (a => 40 , b => 327, p => True ), (a => 41 , b => 326, p => True ), (a => 42 , b => 325, p => True ), (a => 43 , b => 324, p => True ), (a => 44 , b => 323, p => True ), (a => 45 , b => 322, p => True ), (a => 46 , b => 321, p => True ), (a => 47 , b => 320, p => True ), (a => 48 , b => 319, p => True ), (a => 49 , b => 318, p => True ), (a => 50 , b => 317, p => True ), (a => 51 , b => 316, p => True ), (a => 52 , b => 315, p => True ), (a => 53 , b => 314, p => True ), (a => 54 , b => 313, p => True ), (a => 55 , b => 312, p => True ), (a => 56 , b => 311, p => True ), (a => 57 , b => 310, p => True ), (a => 58 , b => 309, p => True ), (a => 59 , b => 308, p => True ), (a => 60 , b => 307, p => True ), (a => 61 , b => 306, p => True ), (a => 62 , b => 305, p => True ), (a => 63 , b => 304, p => True ), (a => 64 , b => 303, p => True ), (a => 65 , b => 302, p => True ), (a => 66 , b => 301, p => True ), (a => 67 , b => 300, p => True ), (a => 68 , b => 299, p => True ), (a => 69 , b => 298, p => True ), (a => 70 , b => 297, p => True ), (a => 71 , b => 296, p => True ), (a => 72 , b => 295, p => True ), (a => 73 , b => 294, p => True ), (a => 74 , b => 293, p => True ), (a => 75 , b => 292, p => True ), (a => 76 , b => 291, p => True ), (a => 77 , b => 290, p => True ), (a => 78 , b => 289, p => True ), (a => 79 , b => 288, p => True ), (a => 80 , b => 287, p => True ), (a => 81 , b => 286, p => True ), (a => 82 , b => 285, p => True ), (a => 83 , b => 284, p => True ), (a => 84 , b => 283, p => True ), (a => 85 , b => 282, p => True ), (a => 86 , b => 281, p => True ), (a => 87 , b => 280, p => True ), (a => 88 , b => 279, p => True ), (a => 89 , b => 278, p => True ), (a => 90 , b => 277, p => True ), (a => 91 , b => 276, p => True ), (a => 92 , b => 275, p => True ), (a => 93 , b => 274, p => True ), (a => 94 , b => 273, p => True ), (a => 95 , b => 272, p => True ), (a => 96 , b => 271, p => True ), (a => 97 , b => 270, p => True ), (a => 98 , b => 269, p => True ), (a => 99 , b => 268, p => True ), (a => 100, b => 267, p => True ), (a => 101, b => 266, p => True ), (a => 102, b => 265, p => True ), (a => 103, b => 264, p => True ), (a => 104, b => 263, p => True ), (a => 105, b => 262, p => True ), (a => 106, b => 261, p => True ), (a => 107, b => 260, p => True ), (a => 108, b => 259, p => True ), (a => 109, b => 258, p => True ), (a => 110, b => 257, p => True ), (a => 111, b => 256, p => True ), (a => 112, b => 255, p => True ), (a => 113, b => 254, p => True ), (a => 114, b => 253, p => True ), (a => 115, b => 252, p => True ), (a => 116, b => 251, p => True ), (a => 117, b => 250, p => True ), (a => 118, b => 249, p => True ), (a => 119, b => 248, p => True ), (a => 120, b => 247, p => True ), (a => 121, b => 246, p => True ), (a => 122, b => 245, p => True ), (a => 123, b => 244, p => True ), (a => 124, b => 243, p => True ), (a => 125, b => 242, p => True ), (a => 126, b => 241, p => True ), (a => 127, b => 240, p => True ), (a => 128, b => 239, p => True ), (a => 129, b => 238, p => True ), (a => 130, b => 237, p => True ), (a => 131, b => 236, p => True ), (a => 132, b => 235, p => True ), (a => 133, b => 234, p => True ), (a => 134, b => 233, p => True ), (a => 135, b => 232, p => True ), (a => 136, b => 231, p => True ), (a => 137, b => 230, p => True ), (a => 138, b => 229, p => True ), (a => 139, b => 228, p => True ), (a => 140, b => 227, p => True ), (a => 141, b => 226, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 146, b => 221, p => True ), (a => 147, b => 220, p => True ), (a => 148, b => 219, p => True ), (a => 149, b => 218, p => True ), (a => 150, b => 217, p => True ), (a => 151, b => 216, p => True ), (a => 152, b => 215, p => True ), (a => 153, b => 214, p => True ), (a => 154, b => 213, p => True ), (a => 155, b => 212, p => True ), (a => 156, b => 211, p => True ), (a => 157, b => 210, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 162, b => 205, p => True ), (a => 163, b => 204, p => True ), (a => 164, b => 203, p => True ), (a => 165, b => 202, p => True ), (a => 166, b => 201, p => True ), (a => 167, b => 200, p => True ), (a => 168, b => 199, p => True ), (a => 169, b => 198, p => True ), (a => 170, b => 197, p => True ), (a => 171, b => 196, p => True ), (a => 172, b => 195, p => True ), (a => 173, b => 194, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True ), (a => 178, b => 189, p => True ), (a => 179, b => 188, p => True ), (a => 180, b => 187, p => True ), (a => 181, b => 186, p => True ), (a => 182, b => 185, p => True ), (a => 183, b => 184, p => True )),
                    ((a => 12 , b => 16 , p => False), (a => 6  , b => 10 , p => False), (a => 14 , b => 18 , p => False), (a => 5  , b => 9  , p => False), (a => 13 , b => 17 , p => False), (a => 7  , b => 11 , p => False), (a => 15 , b => 19 , p => False), (a => 2  , b => 4  , p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 3  , b => 349, p => True ), (a => 8  , b => 348, p => True ), (a => 20 , b => 347, p => True ), (a => 21 , b => 346, p => True ), (a => 22 , b => 345, p => True ), (a => 23 , b => 344, p => True ), (a => 24 , b => 343, p => True ), (a => 25 , b => 342, p => True ), (a => 26 , b => 341, p => True ), (a => 27 , b => 340, p => True ), (a => 28 , b => 339, p => True ), (a => 29 , b => 338, p => True ), (a => 30 , b => 337, p => True ), (a => 31 , b => 336, p => True ), (a => 32 , b => 335, p => True ), (a => 33 , b => 334, p => True ), (a => 34 , b => 333, p => True ), (a => 35 , b => 332, p => True ), (a => 36 , b => 331, p => True ), (a => 37 , b => 330, p => True ), (a => 38 , b => 329, p => True ), (a => 39 , b => 328, p => True ), (a => 40 , b => 327, p => True ), (a => 41 , b => 326, p => True ), (a => 42 , b => 325, p => True ), (a => 43 , b => 324, p => True ), (a => 44 , b => 323, p => True ), (a => 45 , b => 322, p => True ), (a => 46 , b => 321, p => True ), (a => 47 , b => 320, p => True ), (a => 48 , b => 319, p => True ), (a => 49 , b => 318, p => True ), (a => 50 , b => 317, p => True ), (a => 51 , b => 316, p => True ), (a => 52 , b => 315, p => True ), (a => 53 , b => 314, p => True ), (a => 54 , b => 313, p => True ), (a => 55 , b => 312, p => True ), (a => 56 , b => 311, p => True ), (a => 57 , b => 310, p => True ), (a => 58 , b => 309, p => True ), (a => 59 , b => 308, p => True ), (a => 60 , b => 307, p => True ), (a => 61 , b => 306, p => True ), (a => 62 , b => 305, p => True ), (a => 63 , b => 304, p => True ), (a => 64 , b => 303, p => True ), (a => 65 , b => 302, p => True ), (a => 66 , b => 301, p => True ), (a => 67 , b => 300, p => True ), (a => 68 , b => 299, p => True ), (a => 69 , b => 298, p => True ), (a => 70 , b => 297, p => True ), (a => 71 , b => 296, p => True ), (a => 72 , b => 295, p => True ), (a => 73 , b => 294, p => True ), (a => 74 , b => 293, p => True ), (a => 75 , b => 292, p => True ), (a => 76 , b => 291, p => True ), (a => 77 , b => 290, p => True ), (a => 78 , b => 289, p => True ), (a => 79 , b => 288, p => True ), (a => 80 , b => 287, p => True ), (a => 81 , b => 286, p => True ), (a => 82 , b => 285, p => True ), (a => 83 , b => 284, p => True ), (a => 84 , b => 283, p => True ), (a => 85 , b => 282, p => True ), (a => 86 , b => 281, p => True ), (a => 87 , b => 280, p => True ), (a => 88 , b => 279, p => True ), (a => 89 , b => 278, p => True ), (a => 90 , b => 277, p => True ), (a => 91 , b => 276, p => True ), (a => 92 , b => 275, p => True ), (a => 93 , b => 274, p => True ), (a => 94 , b => 273, p => True ), (a => 95 , b => 272, p => True ), (a => 96 , b => 271, p => True ), (a => 97 , b => 270, p => True ), (a => 98 , b => 269, p => True ), (a => 99 , b => 268, p => True ), (a => 100, b => 267, p => True ), (a => 101, b => 266, p => True ), (a => 102, b => 265, p => True ), (a => 103, b => 264, p => True ), (a => 104, b => 263, p => True ), (a => 105, b => 262, p => True ), (a => 106, b => 261, p => True ), (a => 107, b => 260, p => True ), (a => 108, b => 259, p => True ), (a => 109, b => 258, p => True ), (a => 110, b => 257, p => True ), (a => 111, b => 256, p => True ), (a => 112, b => 255, p => True ), (a => 113, b => 254, p => True ), (a => 114, b => 253, p => True ), (a => 115, b => 252, p => True ), (a => 116, b => 251, p => True ), (a => 117, b => 250, p => True ), (a => 118, b => 249, p => True ), (a => 119, b => 248, p => True ), (a => 120, b => 247, p => True ), (a => 121, b => 246, p => True ), (a => 122, b => 245, p => True ), (a => 123, b => 244, p => True ), (a => 124, b => 243, p => True ), (a => 125, b => 242, p => True ), (a => 126, b => 241, p => True ), (a => 127, b => 240, p => True ), (a => 128, b => 239, p => True ), (a => 129, b => 238, p => True ), (a => 130, b => 237, p => True ), (a => 131, b => 236, p => True ), (a => 132, b => 235, p => True ), (a => 133, b => 234, p => True ), (a => 134, b => 233, p => True ), (a => 135, b => 232, p => True ), (a => 136, b => 231, p => True ), (a => 137, b => 230, p => True ), (a => 138, b => 229, p => True ), (a => 139, b => 228, p => True ), (a => 140, b => 227, p => True ), (a => 141, b => 226, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 146, b => 221, p => True ), (a => 147, b => 220, p => True ), (a => 148, b => 219, p => True ), (a => 149, b => 218, p => True ), (a => 150, b => 217, p => True ), (a => 151, b => 216, p => True ), (a => 152, b => 215, p => True ), (a => 153, b => 214, p => True ), (a => 154, b => 213, p => True ), (a => 155, b => 212, p => True ), (a => 156, b => 211, p => True ), (a => 157, b => 210, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 162, b => 205, p => True ), (a => 163, b => 204, p => True ), (a => 164, b => 203, p => True ), (a => 165, b => 202, p => True ), (a => 166, b => 201, p => True ), (a => 167, b => 200, p => True ), (a => 168, b => 199, p => True ), (a => 169, b => 198, p => True ), (a => 170, b => 197, p => True ), (a => 171, b => 196, p => True ), (a => 172, b => 195, p => True ), (a => 173, b => 194, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True ), (a => 178, b => 189, p => True ), (a => 179, b => 188, p => True ), (a => 180, b => 187, p => True ), (a => 181, b => 186, p => True ), (a => 182, b => 185, p => True ), (a => 183, b => 184, p => True )),
                    ((a => 6  , b => 8  , p => False), (a => 10 , b => 12 , p => False), (a => 14 , b => 16 , p => False), (a => 3  , b => 5  , p => False), (a => 7  , b => 9  , p => False), (a => 11 , b => 13 , p => False), (a => 15 , b => 17 , p => False), (a => 1  , b => 2  , p => False), (a => 0  , b => 351, p => True ), (a => 4  , b => 350, p => True ), (a => 18 , b => 349, p => True ), (a => 19 , b => 348, p => True ), (a => 20 , b => 347, p => True ), (a => 21 , b => 346, p => True ), (a => 22 , b => 345, p => True ), (a => 23 , b => 344, p => True ), (a => 24 , b => 343, p => True ), (a => 25 , b => 342, p => True ), (a => 26 , b => 341, p => True ), (a => 27 , b => 340, p => True ), (a => 28 , b => 339, p => True ), (a => 29 , b => 338, p => True ), (a => 30 , b => 337, p => True ), (a => 31 , b => 336, p => True ), (a => 32 , b => 335, p => True ), (a => 33 , b => 334, p => True ), (a => 34 , b => 333, p => True ), (a => 35 , b => 332, p => True ), (a => 36 , b => 331, p => True ), (a => 37 , b => 330, p => True ), (a => 38 , b => 329, p => True ), (a => 39 , b => 328, p => True ), (a => 40 , b => 327, p => True ), (a => 41 , b => 326, p => True ), (a => 42 , b => 325, p => True ), (a => 43 , b => 324, p => True ), (a => 44 , b => 323, p => True ), (a => 45 , b => 322, p => True ), (a => 46 , b => 321, p => True ), (a => 47 , b => 320, p => True ), (a => 48 , b => 319, p => True ), (a => 49 , b => 318, p => True ), (a => 50 , b => 317, p => True ), (a => 51 , b => 316, p => True ), (a => 52 , b => 315, p => True ), (a => 53 , b => 314, p => True ), (a => 54 , b => 313, p => True ), (a => 55 , b => 312, p => True ), (a => 56 , b => 311, p => True ), (a => 57 , b => 310, p => True ), (a => 58 , b => 309, p => True ), (a => 59 , b => 308, p => True ), (a => 60 , b => 307, p => True ), (a => 61 , b => 306, p => True ), (a => 62 , b => 305, p => True ), (a => 63 , b => 304, p => True ), (a => 64 , b => 303, p => True ), (a => 65 , b => 302, p => True ), (a => 66 , b => 301, p => True ), (a => 67 , b => 300, p => True ), (a => 68 , b => 299, p => True ), (a => 69 , b => 298, p => True ), (a => 70 , b => 297, p => True ), (a => 71 , b => 296, p => True ), (a => 72 , b => 295, p => True ), (a => 73 , b => 294, p => True ), (a => 74 , b => 293, p => True ), (a => 75 , b => 292, p => True ), (a => 76 , b => 291, p => True ), (a => 77 , b => 290, p => True ), (a => 78 , b => 289, p => True ), (a => 79 , b => 288, p => True ), (a => 80 , b => 287, p => True ), (a => 81 , b => 286, p => True ), (a => 82 , b => 285, p => True ), (a => 83 , b => 284, p => True ), (a => 84 , b => 283, p => True ), (a => 85 , b => 282, p => True ), (a => 86 , b => 281, p => True ), (a => 87 , b => 280, p => True ), (a => 88 , b => 279, p => True ), (a => 89 , b => 278, p => True ), (a => 90 , b => 277, p => True ), (a => 91 , b => 276, p => True ), (a => 92 , b => 275, p => True ), (a => 93 , b => 274, p => True ), (a => 94 , b => 273, p => True ), (a => 95 , b => 272, p => True ), (a => 96 , b => 271, p => True ), (a => 97 , b => 270, p => True ), (a => 98 , b => 269, p => True ), (a => 99 , b => 268, p => True ), (a => 100, b => 267, p => True ), (a => 101, b => 266, p => True ), (a => 102, b => 265, p => True ), (a => 103, b => 264, p => True ), (a => 104, b => 263, p => True ), (a => 105, b => 262, p => True ), (a => 106, b => 261, p => True ), (a => 107, b => 260, p => True ), (a => 108, b => 259, p => True ), (a => 109, b => 258, p => True ), (a => 110, b => 257, p => True ), (a => 111, b => 256, p => True ), (a => 112, b => 255, p => True ), (a => 113, b => 254, p => True ), (a => 114, b => 253, p => True ), (a => 115, b => 252, p => True ), (a => 116, b => 251, p => True ), (a => 117, b => 250, p => True ), (a => 118, b => 249, p => True ), (a => 119, b => 248, p => True ), (a => 120, b => 247, p => True ), (a => 121, b => 246, p => True ), (a => 122, b => 245, p => True ), (a => 123, b => 244, p => True ), (a => 124, b => 243, p => True ), (a => 125, b => 242, p => True ), (a => 126, b => 241, p => True ), (a => 127, b => 240, p => True ), (a => 128, b => 239, p => True ), (a => 129, b => 238, p => True ), (a => 130, b => 237, p => True ), (a => 131, b => 236, p => True ), (a => 132, b => 235, p => True ), (a => 133, b => 234, p => True ), (a => 134, b => 233, p => True ), (a => 135, b => 232, p => True ), (a => 136, b => 231, p => True ), (a => 137, b => 230, p => True ), (a => 138, b => 229, p => True ), (a => 139, b => 228, p => True ), (a => 140, b => 227, p => True ), (a => 141, b => 226, p => True ), (a => 142, b => 225, p => True ), (a => 143, b => 224, p => True ), (a => 144, b => 223, p => True ), (a => 145, b => 222, p => True ), (a => 146, b => 221, p => True ), (a => 147, b => 220, p => True ), (a => 148, b => 219, p => True ), (a => 149, b => 218, p => True ), (a => 150, b => 217, p => True ), (a => 151, b => 216, p => True ), (a => 152, b => 215, p => True ), (a => 153, b => 214, p => True ), (a => 154, b => 213, p => True ), (a => 155, b => 212, p => True ), (a => 156, b => 211, p => True ), (a => 157, b => 210, p => True ), (a => 158, b => 209, p => True ), (a => 159, b => 208, p => True ), (a => 160, b => 207, p => True ), (a => 161, b => 206, p => True ), (a => 162, b => 205, p => True ), (a => 163, b => 204, p => True ), (a => 164, b => 203, p => True ), (a => 165, b => 202, p => True ), (a => 166, b => 201, p => True ), (a => 167, b => 200, p => True ), (a => 168, b => 199, p => True ), (a => 169, b => 198, p => True ), (a => 170, b => 197, p => True ), (a => 171, b => 196, p => True ), (a => 172, b => 195, p => True ), (a => 173, b => 194, p => True ), (a => 174, b => 193, p => True ), (a => 175, b => 192, p => True ), (a => 176, b => 191, p => True ), (a => 177, b => 190, p => True ), (a => 178, b => 189, p => True ), (a => 179, b => 188, p => True ), (a => 180, b => 187, p => True ), (a => 181, b => 186, p => True ), (a => 182, b => 185, p => True ), (a => 183, b => 184, p => True )),
                    ((a => 3  , b => 4  , p => False), (a => 5  , b => 6  , p => False), (a => 7  , b => 8  , p => False), (a => 9  , b => 10 , p => False), (a => 11 , b => 12 , p => False), (a => 13 , b => 14 , p => False), (a => 15 , b => 16 , p => False), (a => 0  , b => 351, p => True ), (a => 1  , b => 350, p => True ), (a => 2  , b => 349, p => True ), (a => 17 , b => 348, p => True ), (a => 18 , b => 347, p => True ), (a => 19 , b => 346, p => True ), (a => 20 , b => 345, p => True ), (a => 21 , b => 344, p => True ), (a => 22 , b => 343, p => True ), (a => 23 , b => 342, p => True ), (a => 24 , b => 341, p => True ), (a => 25 , b => 340, p => True ), (a => 26 , b => 339, p => True ), (a => 27 , b => 338, p => True ), (a => 28 , b => 337, p => True ), (a => 29 , b => 336, p => True ), (a => 30 , b => 335, p => True ), (a => 31 , b => 334, p => True ), (a => 32 , b => 333, p => True ), (a => 33 , b => 332, p => True ), (a => 34 , b => 331, p => True ), (a => 35 , b => 330, p => True ), (a => 36 , b => 329, p => True ), (a => 37 , b => 328, p => True ), (a => 38 , b => 327, p => True ), (a => 39 , b => 326, p => True ), (a => 40 , b => 325, p => True ), (a => 41 , b => 324, p => True ), (a => 42 , b => 323, p => True ), (a => 43 , b => 322, p => True ), (a => 44 , b => 321, p => True ), (a => 45 , b => 320, p => True ), (a => 46 , b => 319, p => True ), (a => 47 , b => 318, p => True ), (a => 48 , b => 317, p => True ), (a => 49 , b => 316, p => True ), (a => 50 , b => 315, p => True ), (a => 51 , b => 314, p => True ), (a => 52 , b => 313, p => True ), (a => 53 , b => 312, p => True ), (a => 54 , b => 311, p => True ), (a => 55 , b => 310, p => True ), (a => 56 , b => 309, p => True ), (a => 57 , b => 308, p => True ), (a => 58 , b => 307, p => True ), (a => 59 , b => 306, p => True ), (a => 60 , b => 305, p => True ), (a => 61 , b => 304, p => True ), (a => 62 , b => 303, p => True ), (a => 63 , b => 302, p => True ), (a => 64 , b => 301, p => True ), (a => 65 , b => 300, p => True ), (a => 66 , b => 299, p => True ), (a => 67 , b => 298, p => True ), (a => 68 , b => 297, p => True ), (a => 69 , b => 296, p => True ), (a => 70 , b => 295, p => True ), (a => 71 , b => 294, p => True ), (a => 72 , b => 293, p => True ), (a => 73 , b => 292, p => True ), (a => 74 , b => 291, p => True ), (a => 75 , b => 290, p => True ), (a => 76 , b => 289, p => True ), (a => 77 , b => 288, p => True ), (a => 78 , b => 287, p => True ), (a => 79 , b => 286, p => True ), (a => 80 , b => 285, p => True ), (a => 81 , b => 284, p => True ), (a => 82 , b => 283, p => True ), (a => 83 , b => 282, p => True ), (a => 84 , b => 281, p => True ), (a => 85 , b => 280, p => True ), (a => 86 , b => 279, p => True ), (a => 87 , b => 278, p => True ), (a => 88 , b => 277, p => True ), (a => 89 , b => 276, p => True ), (a => 90 , b => 275, p => True ), (a => 91 , b => 274, p => True ), (a => 92 , b => 273, p => True ), (a => 93 , b => 272, p => True ), (a => 94 , b => 271, p => True ), (a => 95 , b => 270, p => True ), (a => 96 , b => 269, p => True ), (a => 97 , b => 268, p => True ), (a => 98 , b => 267, p => True ), (a => 99 , b => 266, p => True ), (a => 100, b => 265, p => True ), (a => 101, b => 264, p => True ), (a => 102, b => 263, p => True ), (a => 103, b => 262, p => True ), (a => 104, b => 261, p => True ), (a => 105, b => 260, p => True ), (a => 106, b => 259, p => True ), (a => 107, b => 258, p => True ), (a => 108, b => 257, p => True ), (a => 109, b => 256, p => True ), (a => 110, b => 255, p => True ), (a => 111, b => 254, p => True ), (a => 112, b => 253, p => True ), (a => 113, b => 252, p => True ), (a => 114, b => 251, p => True ), (a => 115, b => 250, p => True ), (a => 116, b => 249, p => True ), (a => 117, b => 248, p => True ), (a => 118, b => 247, p => True ), (a => 119, b => 246, p => True ), (a => 120, b => 245, p => True ), (a => 121, b => 244, p => True ), (a => 122, b => 243, p => True ), (a => 123, b => 242, p => True ), (a => 124, b => 241, p => True ), (a => 125, b => 240, p => True ), (a => 126, b => 239, p => True ), (a => 127, b => 238, p => True ), (a => 128, b => 237, p => True ), (a => 129, b => 236, p => True ), (a => 130, b => 235, p => True ), (a => 131, b => 234, p => True ), (a => 132, b => 233, p => True ), (a => 133, b => 232, p => True ), (a => 134, b => 231, p => True ), (a => 135, b => 230, p => True ), (a => 136, b => 229, p => True ), (a => 137, b => 228, p => True ), (a => 138, b => 227, p => True ), (a => 139, b => 226, p => True ), (a => 140, b => 225, p => True ), (a => 141, b => 224, p => True ), (a => 142, b => 223, p => True ), (a => 143, b => 222, p => True ), (a => 144, b => 221, p => True ), (a => 145, b => 220, p => True ), (a => 146, b => 219, p => True ), (a => 147, b => 218, p => True ), (a => 148, b => 217, p => True ), (a => 149, b => 216, p => True ), (a => 150, b => 215, p => True ), (a => 151, b => 214, p => True ), (a => 152, b => 213, p => True ), (a => 153, b => 212, p => True ), (a => 154, b => 211, p => True ), (a => 155, b => 210, p => True ), (a => 156, b => 209, p => True ), (a => 157, b => 208, p => True ), (a => 158, b => 207, p => True ), (a => 159, b => 206, p => True ), (a => 160, b => 205, p => True ), (a => 161, b => 204, p => True ), (a => 162, b => 203, p => True ), (a => 163, b => 202, p => True ), (a => 164, b => 201, p => True ), (a => 165, b => 200, p => True ), (a => 166, b => 199, p => True ), (a => 167, b => 198, p => True ), (a => 168, b => 197, p => True ), (a => 169, b => 196, p => True ), (a => 170, b => 195, p => True ), (a => 171, b => 194, p => True ), (a => 172, b => 193, p => True ), (a => 173, b => 192, p => True ), (a => 174, b => 191, p => True ), (a => 175, b => 190, p => True ), (a => 176, b => 189, p => True ), (a => 177, b => 188, p => True ), (a => 178, b => 187, p => True ), (a => 179, b => 186, p => True ), (a => 180, b => 185, p => True ), (a => 181, b => 184, p => True ), (a => 182, b => 183, p => True ))
                    );
					

			when others => return empty_cfg;

		end case;
	end function get_cfg;


	function get_stg(I : integer; D: integer) return stages_a is
        begin
            case I is
                when 64  =>
                    case D is
                        when 4 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20|;
                        return    ( False, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True);
                        -- total number of registered stages: 4.
                        when 5 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20|;
                        return    ( False, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 5.
                        when 6 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20|;
                        return    ( False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 6.
                        when 7 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20|;
                        return    ( False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True);
                        -- total number of registered stages: 7.
                        when 8 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20|;
                        return    ( False,  True, False, False,  True, False,  True, False, False,  True, False, False,  True, False,  True, False, False,  True, False, False,  True);
                        -- total number of registered stages: 8.
                        when 9 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20|;
                        return    ( False, False,  True, False,  True, False, False,  True, False,  True, False,  True, False, False,  True, False,  True, False,  True, False,  True);
                        -- total number of registered stages: 9.
                        when others =>
                        null;
                     end case;

                when 88  =>
                    case D is
                        when 4 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27|;
                        return    ( False, False, False, False, False, False,  True, False, False, False, False, False, False,  True, False, False, False, False, False, False,  True, False, False, False, False, False, False,  True);
                        -- total number of registered stages: 4.
                        when 5 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27|;
                        return    ( False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False, False,  True);
                        -- total number of registered stages: 5.
                        when 6 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27|;
                        return    ( False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True);
                        -- total number of registered stages: 6.
                        when 7 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27|;
                        return    ( False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 7.
                        when 8 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27|;
                        return    ( False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 8.
                        when 9 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27|;
                        return    ( False, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True);
                        -- total number of registered stages: 9.
                        when others =>
                                                null;
                    end case;
                when 352 =>
                    case D is
                        when 6 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False, False, False, False, False,  True, False, False, False, False, False, False,  True, False, False, False, False, False, False, False,  True, False, False, False, False, False, False,  True, False, False, False, False, False, False,  True, False, False, False, False, False, False,  True);
                        -- total number of registered stages: 6.
                        when 7 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False, False,  True);
                        -- total number of registered stages: 7.
                        when 8 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False, False,  True);
                        -- total number of registered stages: 8.
                        when 9 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True, False, False, False, False,  True);
                        -- total number of registered stages: 9.
                        when 10 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False, False,  True, False, False, False,  True, False, False, False, False,  True, False, False, False,  True, False, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False, False,  True, False, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 10.
                        when 11 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 11.
                        when 12 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False,  True, False, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False, False,  True);
                        -- total number of registered stages: 12.
                        when 13 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False,  True);
                        -- total number of registered stages: 13.
                        when 14 =>
                        -- Registered stages configuration
                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31,    32,    33,    34,    35,    36,    37,    38,    39,    40,    41,    42,    43|;
                        return    ( False, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True, False, False,  True);
                        -- total number of registered stages: 14.

                    when others =>
                        null;
                    end case;

                when others => return (False, False);

            end case;
        end function get_stg;


	function to_array(data : std_logic_vector; N : integer) return muon_a is
		variable muon : muon_a(0 to N - 1);
	begin
		for i in muon'range loop
			muon(i).pt  := data((i + 1) * word_w - 1 - IDX_WIDTH downto i * word_w);
			muon(i).idx := data((i + 1) * word_w - 1 downto i * word_w + PT_WIDTH);
		end loop;
		return muon;
	end to_array;
	
	function to_sel_array(data : std_logic_vector; N : integer) return muon_sel_a is
		variable muon : muon_sel_a(0 to N - 1);
	begin
		for i in muon'range loop
			muon(i).pt  := data((i + 1) * PT_WIDTH - 1 downto i * PT_WIDTH);			
		end loop;
		return muon;
	end to_sel_array;

	function to_stdv(muon : muon_a; N : integer) return std_logic_vector is
		variable vector : std_logic_vector(N * word_w - 1 downto 0);
	begin
		for i in muon'range loop
			vector((i + 1) * word_w - 1 - IDX_WIDTH downto i * word_w) := muon(i).pt;
			vector((i + 1) * word_w - 1 downto i * word_w + PT_WIDTH)  := muon(i).idx;
		end loop;
		return vector;
	end to_stdv;

end package body csn_pkg;
