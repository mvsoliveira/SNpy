library ieee;
use ieee.std_logic_1164.all;
use IEEE.math_real.all;

package csn_pkg is

  constant MUON_NUMBER : integer := 352;
  constant IDX_WIDTH   : integer := integer(ceil(log(real(MUON_NUMBER), real(2))));
  constant PT_WIDTH    : integer := 4;
  constant ROI_WIDTH   : integer := 8;
  constant FLAGS_WIDTH : integer := 4;
  constant in_word_w   : integer := PT_WIDTH + ROI_WIDTH + FLAGS_WIDTH;
  constant out_word_w  : integer := PT_WIDTH + ROI_WIDTH + FLAGS_WIDTH + IDX_WIDTH;

  type muon_type is record
    idx   : std_logic_vector(IDX_WIDTH - 1 downto 0);
    pt    : std_logic_vector(PT_WIDTH - 1 downto 0);
    roi   : std_logic_vector(ROI_WIDTH - 1 downto 0);
    flags : std_logic_vector(FLAGS_WIDTH - 1 downto 0);
  end record;

  type muon_sort_type is record
    pt  : std_logic_vector(PT_WIDTH - 1 downto 0);
    idx : std_logic_vector(IDX_WIDTH - 1 downto 0);
  end record;

  type muon_a is array (natural range <>) of muon_type;
  type muon_sort_a is array (natural range <>) of muon_sort_type;

  type cmp_cfg is record
    a : natural;
    b : natural;
    p : boolean;
  end record;

  -- has to be array of array instead of (x,y) array because of issues with synplify
  type pair_cmp_cfg is array (natural range <>) of cmp_cfg;
  type cfg_net_t is array (natural range <>) of pair_cmp_cfg;
  type stages_a is array (natural range <>) of boolean;

  function to_array(data : std_logic_vector; N : integer) return muon_a;
  function to_stdv(muon  : muon_a; N : integer) return std_logic_vector;

  --type cfg_net_t is array (natural range <>, natural range <>) of cmp_cfg;
  function get_cfg(I         : integer) return cfg_net_t;
  function get_stg(I         : integer; D : integer) return stages_a;
  function get_stg_off(depth : integer; D : integer; Off : integer) return stages_a;

  constant empty_cfg : cfg_net_t := (
    ((a => 0, b => 1, p => false), (a => 2, b => 3, p => false)),
    ((a => 0, b => 2, p => false), (a => 1, b => 3, p => false)),
    ((a => 1, b => 2, p => false), (a => 0, b => 3, p => true))
    );

end package csn_pkg;

package body csn_pkg is

  function get_cfg(I : integer) return cfg_net_t is
  begin
    case I is
      -- Sherenaz W. Al-Haj Baddar 22-key 12-step SORTING network
      when 22 => return (
        ((a   => 20, b => 21, p => false), (a => 18, b => 19, p => false), (a => 16, b => 17, p => false), (a => 14, b => 15, p => false), (a => 12, b => 13, p => false), (a => 10, b => 11, p => false), (a => 8, b => 9, p => false), (a => 6, b => 7, p => false), (a => 4, b => 5, p => false), (a => 2, b => 3, p => false), (a => 0, b => 1, p => false)),
        ((a   => 17, b => 19, p => false), (a => 13, b => 15, p => false), (a => 9, b => 11, p => false), (a => 5, b => 7, p => false), (a => 1, b => 3, p => false), (a => 18, b => 20, p => false), (a => 12, b => 14, p => false), (a => 8, b => 10, p => false), (a => 4, b => 6, p => false), (a => 0, b => 2, p => false), (a => 16, b => 21, p => false)),
        ((a   => 11, b => 15, p => false), (a => 3, b => 7, p => false), (a => 16, b => 18, p => false), (a => 19, b => 21, p => false), (a => 10, b => 14, p => false), (a => 2, b => 6, p => false), (a => 17, b => 20, p => false), (a => 9, b => 13, p => false), (a => 1, b => 5, p => false), (a => 8, b => 12, p => false), (a => 0, b => 4, p => false)),
        ((a   => 4, b => 12, p => false), (a => 17, b => 19, p => false), (a => 6, b => 14, p => false), (a => 2, b => 10, p => false), (a => 11, b => 21, p => false), (a => 5, b => 13, p => false), (a => 9, b => 18, p => false), (a => 0, b => 8, p => false), (a => 3, b => 20, p => false), (a => 1, b => 16, p => false), (a => 7, b => 15, p => false)),
        ((a   => 14, b => 21, p => false), (a => 1, b => 4, p => false), (a => 7, b => 8, p => false), (a => 6, b => 18, p => false), (a => 3, b => 12, p => false), (a => 13, b => 20, p => false), (a => 10, b => 19, p => false), (a => 2, b => 9, p => false), (a => 5, b => 17, p => false), (a => 11, b => 16, p => false), (a => 0, b => 15, p => true)),
        ((a   => 0, b => 1, p => false), (a => 15, b => 21, p => false), (a => 3, b => 9, p => false), (a => 13, b => 18, p => false), (a => 5, b => 7, p => false), (a => 8, b => 19, p => false), (a => 12, b => 16, p => false), (a => 6, b => 11, p => false), (a => 14, b => 17, p => false), (a => 4, b => 10, p => false), (a => 2, b => 20, p => true)),
        ((a   => 1, b => 5, p => false), (a => 7, b => 9, p => false), (a => 10, b => 11, p => false), (a => 12, b => 14, p => false), (a => 16, b => 17, p => false), (a => 18, b => 20, p => false), (a => 2, b => 3, p => false), (a => 4, b => 6, p => false), (a => 8, b => 13, p => false), (a => 15, b => 19, p => false), (a => 0, b => 21, p => true)),
        ((a   => 1, b => 2, p => false), (a => 4, b => 5, p => false), (a => 7, b => 10, p => false), (a => 13, b => 14, p => false), (a => 16, b => 18, p => false), (a => 19, b => 20, p => false), (a => 3, b => 6, p => false), (a => 8, b => 12, p => false), (a => 15, b => 17, p => false), (a => 9, b => 11, p => false), (a => 0, b => 21, p => true)),
        ((a   => 2, b => 3, p => false), (a => 5, b => 7, p => false), (a => 9, b => 10, p => false), (a => 12, b => 13, p => false), (a => 14, b => 15, p => false), (a => 18, b => 19, p => false), (a => 6, b => 8, p => false), (a => 11, b => 16, p => false), (a => 0, b => 21, p => true), (a => 1, b => 20, p => true), (a => 4, b => 17, p => true)),
        ((a   => 2, b => 4, p => false), (a => 6, b => 7, p => false), (a => 8, b => 9, p => false), (a => 10, b => 12, p => false), (a => 14, b => 16, p => false), (a => 3, b => 5, p => false), (a => 11, b => 13, p => false), (a => 15, b => 18, p => false), (a => 0, b => 21, p => true), (a => 1, b => 20, p => true), (a => 17, b => 19, p => true)),
        ((a   => 3, b => 4, p => false), (a => 5, b => 6, p => false), (a => 7, b => 8, p => false), (a => 9, b => 10, p => false), (a => 11, b => 12, p => false), (a => 13, b => 14, p => false), (a => 15, b => 16, p => false), (a => 0, b => 21, p => true), (a => 1, b => 20, p => true), (a => 2, b => 19, p => true), (a => 17, b => 18, p => true)),
        ((a   => 4, b => 5, p => false), (a => 6, b => 7, p => false), (a => 8, b => 9, p => false), (a => 10, b => 11, p => false), (a => 12, b => 13, p => false), (a => 14, b => 15, p => false), (a => 0, b => 21, p => true), (a => 1, b => 20, p => true), (a => 2, b => 19, p => true), (a => 3, b => 18, p => true), (a => 16, b => 17, p => true))
        );
      -- M=16,N=16 Batcher Odd-even MERGING network, the two 16-key input sequences have to be sorted 
      when 32 => return (
        ((a   => 0, b => 16, p => false), (a => 8, b => 24, p => false), (a => 4, b => 20, p => false), (a => 12, b => 28, p => false), (a => 2, b => 18, p => false), (a => 10, b => 26, p => false), (a => 6, b => 22, p => false), (a => 14, b => 30, p => false), (a => 1, b => 17, p => false), (a => 9, b => 25, p => false), (a => 5, b => 21, p => false), (a => 13, b => 29, p => false), (a => 3, b => 19, p => false), (a => 11, b => 27, p => false), (a => 7, b => 23, p => false), (a => 15, b => 31, p => false)),
        ((a   => 8, b => 16, p => false), (a => 12, b => 20, p => false), (a => 10, b => 18, p => false), (a => 14, b => 22, p => false), (a => 9, b => 17, p => false), (a => 13, b => 21, p => false), (a => 11, b => 19, p => false), (a => 15, b => 23, p => false), (a => 0, b => 31, p => true), (a => 1, b => 30, p => true), (a => 2, b => 29, p => true), (a => 3, b => 28, p => true), (a => 4, b => 27, p => true), (a => 5, b => 26, p => true), (a => 6, b => 25, p => true), (a => 7, b => 24, p => true)),
        ((a   => 4, b => 8, p => false), (a => 12, b => 16, p => false), (a => 6, b => 10, p => false), (a => 14, b => 18, p => false), (a => 5, b => 9, p => false), (a => 13, b => 17, p => false), (a => 7, b => 11, p => false), (a => 15, b => 19, p => false), (a => 0, b => 31, p => true), (a => 1, b => 30, p => true), (a => 2, b => 29, p => true), (a => 3, b => 28, p => true), (a => 20, b => 27, p => true), (a => 21, b => 26, p => true), (a => 22, b => 25, p => true), (a => 23, b => 24, p => true)),
        ((a   => 2, b => 4, p => false), (a => 6, b => 8, p => false), (a => 10, b => 12, p => false), (a => 14, b => 16, p => false), (a => 3, b => 5, p => false), (a => 7, b => 9, p => false), (a => 11, b => 13, p => false), (a => 15, b => 17, p => false), (a => 0, b => 31, p => true), (a => 1, b => 30, p => true), (a => 18, b => 29, p => true), (a => 19, b => 28, p => true), (a => 20, b => 27, p => true), (a => 21, b => 26, p => true), (a => 22, b => 25, p => true), (a => 23, b => 24, p => true)),
        ((a   => 1, b => 2, p => false), (a => 3, b => 4, p => false), (a => 5, b => 6, p => false), (a => 7, b => 8, p => false), (a => 9, b => 10, p => false), (a => 11, b => 12, p => false), (a => 13, b => 14, p => false), (a => 15, b => 16, p => false), (a => 0, b => 31, p => true), (a => 17, b => 30, p => true), (a => 18, b => 29, p => true), (a => 19, b => 28, p => true), (a => 20, b => 27, p => true), (a => 21, b => 26, p => true), (a => 22, b => 25, p => true), (a => 23, b => 24, p => true))
        );

      when 352 => return (
        ((a    => 20, b => 21, p => false), (a => 42, b => 43, p => false), (a => 64, b => 65, p => false), (a => 86, b => 87, p => false), (a => 108, b => 109, p => false), (a => 130, b => 131, p => false), (a => 152, b => 153, p => false), (a => 174, b => 175, p => false), (a => 196, b => 197, p => false), (a => 218, b => 219, p => false), (a => 240, b => 241, p => false), (a => 262, b => 263, p => false), (a => 284, b => 285, p => false), (a => 306, b => 307, p => false), (a => 328, b => 329, p => false), (a => 350, b => 351, p => false), (a => 18, b => 19, p => false), (a => 40, b => 41, p => false), (a => 62, b => 63, p => false), (a => 84, b => 85, p => false), (a => 106, b => 107, p => false), (a => 128, b => 129, p => false), (a => 150, b => 151, p => false), (a => 172, b => 173, p => false), (a => 194, b => 195, p => false), (a => 216, b => 217, p => false), (a => 238, b => 239, p => false), (a => 260, b => 261, p => false), (a => 282, b => 283, p => false), (a => 304, b => 305, p => false), (a => 326, b => 327, p => false), (a => 348, b => 349, p => false), (a => 16, b => 17, p => false), (a => 38, b => 39, p => false), (a => 60, b => 61, p => false), (a => 82, b => 83, p => false), (a => 104, b => 105, p => false), (a => 126, b => 127, p => false), (a => 148, b => 149, p => false), (a => 170, b => 171, p => false), (a => 192, b => 193, p => false), (a => 214, b => 215, p => false), (a => 236, b => 237, p => false), (a => 258, b => 259, p => false), (a => 280, b => 281, p => false), (a => 302, b => 303, p => false), (a => 324, b => 325, p => false), (a => 346, b => 347, p => false), (a => 14, b => 15, p => false), (a => 36, b => 37, p => false), (a => 58, b => 59, p => false), (a => 80, b => 81, p => false), (a => 102, b => 103, p => false), (a => 124, b => 125, p => false), (a => 146, b => 147, p => false), (a => 168, b => 169, p => false), (a => 190, b => 191, p => false), (a => 212, b => 213, p => false), (a => 234, b => 235, p => false), (a => 256, b => 257, p => false), (a => 278, b => 279, p => false), (a => 300, b => 301, p => false), (a => 322, b => 323, p => false), (a => 344, b => 345, p => false), (a => 12, b => 13, p => false), (a => 34, b => 35, p => false), (a => 56, b => 57, p => false), (a => 78, b => 79, p => false), (a => 100, b => 101, p => false), (a => 122, b => 123, p => false), (a => 144, b => 145, p => false), (a => 166, b => 167, p => false), (a => 188, b => 189, p => false), (a => 210, b => 211, p => false), (a => 232, b => 233, p => false), (a => 254, b => 255, p => false), (a => 276, b => 277, p => false), (a => 298, b => 299, p => false), (a => 320, b => 321, p => false), (a => 342, b => 343, p => false), (a => 10, b => 11, p => false), (a => 32, b => 33, p => false), (a => 54, b => 55, p => false), (a => 76, b => 77, p => false), (a => 98, b => 99, p => false), (a => 120, b => 121, p => false), (a => 142, b => 143, p => false), (a => 164, b => 165, p => false), (a => 186, b => 187, p => false), (a => 208, b => 209, p => false), (a => 230, b => 231, p => false), (a => 252, b => 253, p => false), (a => 274, b => 275, p => false), (a => 296, b => 297, p => false), (a => 318, b => 319, p => false), (a => 340, b => 341, p => false), (a => 8, b => 9, p => false), (a => 30, b => 31, p => false), (a => 52, b => 53, p => false), (a => 74, b => 75, p => false), (a => 96, b => 97, p => false), (a => 118, b => 119, p => false), (a => 140, b => 141, p => false), (a => 162, b => 163, p => false), (a => 184, b => 185, p => false), (a => 206, b => 207, p => false), (a => 228, b => 229, p => false), (a => 250, b => 251, p => false), (a => 272, b => 273, p => false), (a => 294, b => 295, p => false), (a => 316, b => 317, p => false), (a => 338, b => 339, p => false), (a => 6, b => 7, p => false), (a => 28, b => 29, p => false), (a => 50, b => 51, p => false), (a => 72, b => 73, p => false), (a => 94, b => 95, p => false), (a => 116, b => 117, p => false), (a => 138, b => 139, p => false), (a => 160, b => 161, p => false), (a => 182, b => 183, p => false), (a => 204, b => 205, p => false), (a => 226, b => 227, p => false), (a => 248, b => 249, p => false), (a => 270, b => 271, p => false), (a => 292, b => 293, p => false), (a => 314, b => 315, p => false), (a => 336, b => 337, p => false), (a => 4, b => 5, p => false), (a => 26, b => 27, p => false), (a => 48, b => 49, p => false), (a => 70, b => 71, p => false), (a => 92, b => 93, p => false), (a => 114, b => 115, p => false), (a => 136, b => 137, p => false), (a => 158, b => 159, p => false), (a => 180, b => 181, p => false), (a => 202, b => 203, p => false), (a => 224, b => 225, p => false), (a => 246, b => 247, p => false), (a => 268, b => 269, p => false), (a => 290, b => 291, p => false), (a => 312, b => 313, p => false), (a => 334, b => 335, p => false), (a => 2, b => 3, p => false), (a => 24, b => 25, p => false), (a => 46, b => 47, p => false), (a => 68, b => 69, p => false), (a => 90, b => 91, p => false), (a => 112, b => 113, p => false), (a => 134, b => 135, p => false), (a => 156, b => 157, p => false), (a => 178, b => 179, p => false), (a => 200, b => 201, p => false), (a => 222, b => 223, p => false), (a => 244, b => 245, p => false), (a => 266, b => 267, p => false), (a => 288, b => 289, p => false), (a => 310, b => 311, p => false), (a => 332, b => 333, p => false), (a => 0, b => 1, p => false), (a => 22, b => 23, p => false), (a => 44, b => 45, p => false), (a => 66, b => 67, p => false), (a => 88, b => 89, p => false), (a => 110, b => 111, p => false), (a => 132, b => 133, p => false), (a => 154, b => 155, p => false), (a => 176, b => 177, p => false), (a => 198, b => 199, p => false), (a => 220, b => 221, p => false), (a => 242, b => 243, p => false), (a => 264, b => 265, p => false), (a => 286, b => 287, p => false), (a => 308, b => 309, p => false), (a => 330, b => 331, p => false)),
        ((a    => 17, b => 19, p => false), (a => 39, b => 41, p => false), (a => 61, b => 63, p => false), (a => 83, b => 85, p => false), (a => 105, b => 107, p => false), (a => 127, b => 129, p => false), (a => 149, b => 151, p => false), (a => 171, b => 173, p => false), (a => 193, b => 195, p => false), (a => 215, b => 217, p => false), (a => 237, b => 239, p => false), (a => 259, b => 261, p => false), (a => 281, b => 283, p => false), (a => 303, b => 305, p => false), (a => 325, b => 327, p => false), (a => 347, b => 349, p => false), (a => 13, b => 15, p => false), (a => 35, b => 37, p => false), (a => 57, b => 59, p => false), (a => 79, b => 81, p => false), (a => 101, b => 103, p => false), (a => 123, b => 125, p => false), (a => 145, b => 147, p => false), (a => 167, b => 169, p => false), (a => 189, b => 191, p => false), (a => 211, b => 213, p => false), (a => 233, b => 235, p => false), (a => 255, b => 257, p => false), (a => 277, b => 279, p => false), (a => 299, b => 301, p => false), (a => 321, b => 323, p => false), (a => 343, b => 345, p => false), (a => 9, b => 11, p => false), (a => 31, b => 33, p => false), (a => 53, b => 55, p => false), (a => 75, b => 77, p => false), (a => 97, b => 99, p => false), (a => 119, b => 121, p => false), (a => 141, b => 143, p => false), (a => 163, b => 165, p => false), (a => 185, b => 187, p => false), (a => 207, b => 209, p => false), (a => 229, b => 231, p => false), (a => 251, b => 253, p => false), (a => 273, b => 275, p => false), (a => 295, b => 297, p => false), (a => 317, b => 319, p => false), (a => 339, b => 341, p => false), (a => 5, b => 7, p => false), (a => 27, b => 29, p => false), (a => 49, b => 51, p => false), (a => 71, b => 73, p => false), (a => 93, b => 95, p => false), (a => 115, b => 117, p => false), (a => 137, b => 139, p => false), (a => 159, b => 161, p => false), (a => 181, b => 183, p => false), (a => 203, b => 205, p => false), (a => 225, b => 227, p => false), (a => 247, b => 249, p => false), (a => 269, b => 271, p => false), (a => 291, b => 293, p => false), (a => 313, b => 315, p => false), (a => 335, b => 337, p => false), (a => 1, b => 3, p => false), (a => 23, b => 25, p => false), (a => 45, b => 47, p => false), (a => 67, b => 69, p => false), (a => 89, b => 91, p => false), (a => 111, b => 113, p => false), (a => 133, b => 135, p => false), (a => 155, b => 157, p => false), (a => 177, b => 179, p => false), (a => 199, b => 201, p => false), (a => 221, b => 223, p => false), (a => 243, b => 245, p => false), (a => 265, b => 267, p => false), (a => 287, b => 289, p => false), (a => 309, b => 311, p => false), (a => 331, b => 333, p => false), (a => 18, b => 20, p => false), (a => 40, b => 42, p => false), (a => 62, b => 64, p => false), (a => 84, b => 86, p => false), (a => 106, b => 108, p => false), (a => 128, b => 130, p => false), (a => 150, b => 152, p => false), (a => 172, b => 174, p => false), (a => 194, b => 196, p => false), (a => 216, b => 218, p => false), (a => 238, b => 240, p => false), (a => 260, b => 262, p => false), (a => 282, b => 284, p => false), (a => 304, b => 306, p => false), (a => 326, b => 328, p => false), (a => 348, b => 350, p => false), (a => 12, b => 14, p => false), (a => 34, b => 36, p => false), (a => 56, b => 58, p => false), (a => 78, b => 80, p => false), (a => 100, b => 102, p => false), (a => 122, b => 124, p => false), (a => 144, b => 146, p => false), (a => 166, b => 168, p => false), (a => 188, b => 190, p => false), (a => 210, b => 212, p => false), (a => 232, b => 234, p => false), (a => 254, b => 256, p => false), (a => 276, b => 278, p => false), (a => 298, b => 300, p => false), (a => 320, b => 322, p => false), (a => 342, b => 344, p => false), (a => 8, b => 10, p => false), (a => 30, b => 32, p => false), (a => 52, b => 54, p => false), (a => 74, b => 76, p => false), (a => 96, b => 98, p => false), (a => 118, b => 120, p => false), (a => 140, b => 142, p => false), (a => 162, b => 164, p => false), (a => 184, b => 186, p => false), (a => 206, b => 208, p => false), (a => 228, b => 230, p => false), (a => 250, b => 252, p => false), (a => 272, b => 274, p => false), (a => 294, b => 296, p => false), (a => 316, b => 318, p => false), (a => 338, b => 340, p => false), (a => 4, b => 6, p => false), (a => 26, b => 28, p => false), (a => 48, b => 50, p => false), (a => 70, b => 72, p => false), (a => 92, b => 94, p => false), (a => 114, b => 116, p => false), (a => 136, b => 138, p => false), (a => 158, b => 160, p => false), (a => 180, b => 182, p => false), (a => 202, b => 204, p => false), (a => 224, b => 226, p => false), (a => 246, b => 248, p => false), (a => 268, b => 270, p => false), (a => 290, b => 292, p => false), (a => 312, b => 314, p => false), (a => 334, b => 336, p => false), (a => 0, b => 2, p => false), (a => 22, b => 24, p => false), (a => 44, b => 46, p => false), (a => 66, b => 68, p => false), (a => 88, b => 90, p => false), (a => 110, b => 112, p => false), (a => 132, b => 134, p => false), (a => 154, b => 156, p => false), (a => 176, b => 178, p => false), (a => 198, b => 200, p => false), (a => 220, b => 222, p => false), (a => 242, b => 244, p => false), (a => 264, b => 266, p => false), (a => 286, b => 288, p => false), (a => 308, b => 310, p => false), (a => 330, b => 332, p => false), (a => 16, b => 21, p => false), (a => 38, b => 43, p => false), (a => 60, b => 65, p => false), (a => 82, b => 87, p => false), (a => 104, b => 109, p => false), (a => 126, b => 131, p => false), (a => 148, b => 153, p => false), (a => 170, b => 175, p => false), (a => 192, b => 197, p => false), (a => 214, b => 219, p => false), (a => 236, b => 241, p => false), (a => 258, b => 263, p => false), (a => 280, b => 285, p => false), (a => 302, b => 307, p => false), (a => 324, b => 329, p => false), (a => 346, b => 351, p => false)),
        ((a    => 11, b => 15, p => false), (a => 33, b => 37, p => false), (a => 55, b => 59, p => false), (a => 77, b => 81, p => false), (a => 99, b => 103, p => false), (a => 121, b => 125, p => false), (a => 143, b => 147, p => false), (a => 165, b => 169, p => false), (a => 187, b => 191, p => false), (a => 209, b => 213, p => false), (a => 231, b => 235, p => false), (a => 253, b => 257, p => false), (a => 275, b => 279, p => false), (a => 297, b => 301, p => false), (a => 319, b => 323, p => false), (a => 341, b => 345, p => false), (a => 3, b => 7, p => false), (a => 25, b => 29, p => false), (a => 47, b => 51, p => false), (a => 69, b => 73, p => false), (a => 91, b => 95, p => false), (a => 113, b => 117, p => false), (a => 135, b => 139, p => false), (a => 157, b => 161, p => false), (a => 179, b => 183, p => false), (a => 201, b => 205, p => false), (a => 223, b => 227, p => false), (a => 245, b => 249, p => false), (a => 267, b => 271, p => false), (a => 289, b => 293, p => false), (a => 311, b => 315, p => false), (a => 333, b => 337, p => false), (a => 16, b => 18, p => false), (a => 38, b => 40, p => false), (a => 60, b => 62, p => false), (a => 82, b => 84, p => false), (a => 104, b => 106, p => false), (a => 126, b => 128, p => false), (a => 148, b => 150, p => false), (a => 170, b => 172, p => false), (a => 192, b => 194, p => false), (a => 214, b => 216, p => false), (a => 236, b => 238, p => false), (a => 258, b => 260, p => false), (a => 280, b => 282, p => false), (a => 302, b => 304, p => false), (a => 324, b => 326, p => false), (a => 346, b => 348, p => false), (a => 19, b => 21, p => false), (a => 41, b => 43, p => false), (a => 63, b => 65, p => false), (a => 85, b => 87, p => false), (a => 107, b => 109, p => false), (a => 129, b => 131, p => false), (a => 151, b => 153, p => false), (a => 173, b => 175, p => false), (a => 195, b => 197, p => false), (a => 217, b => 219, p => false), (a => 239, b => 241, p => false), (a => 261, b => 263, p => false), (a => 283, b => 285, p => false), (a => 305, b => 307, p => false), (a => 327, b => 329, p => false), (a => 349, b => 351, p => false), (a => 10, b => 14, p => false), (a => 32, b => 36, p => false), (a => 54, b => 58, p => false), (a => 76, b => 80, p => false), (a => 98, b => 102, p => false), (a => 120, b => 124, p => false), (a => 142, b => 146, p => false), (a => 164, b => 168, p => false), (a => 186, b => 190, p => false), (a => 208, b => 212, p => false), (a => 230, b => 234, p => false), (a => 252, b => 256, p => false), (a => 274, b => 278, p => false), (a => 296, b => 300, p => false), (a => 318, b => 322, p => false), (a => 340, b => 344, p => false), (a => 2, b => 6, p => false), (a => 24, b => 28, p => false), (a => 46, b => 50, p => false), (a => 68, b => 72, p => false), (a => 90, b => 94, p => false), (a => 112, b => 116, p => false), (a => 134, b => 138, p => false), (a => 156, b => 160, p => false), (a => 178, b => 182, p => false), (a => 200, b => 204, p => false), (a => 222, b => 226, p => false), (a => 244, b => 248, p => false), (a => 266, b => 270, p => false), (a => 288, b => 292, p => false), (a => 310, b => 314, p => false), (a => 332, b => 336, p => false), (a => 17, b => 20, p => false), (a => 39, b => 42, p => false), (a => 61, b => 64, p => false), (a => 83, b => 86, p => false), (a => 105, b => 108, p => false), (a => 127, b => 130, p => false), (a => 149, b => 152, p => false), (a => 171, b => 174, p => false), (a => 193, b => 196, p => false), (a => 215, b => 218, p => false), (a => 237, b => 240, p => false), (a => 259, b => 262, p => false), (a => 281, b => 284, p => false), (a => 303, b => 306, p => false), (a => 325, b => 328, p => false), (a => 347, b => 350, p => false), (a => 9, b => 13, p => false), (a => 31, b => 35, p => false), (a => 53, b => 57, p => false), (a => 75, b => 79, p => false), (a => 97, b => 101, p => false), (a => 119, b => 123, p => false), (a => 141, b => 145, p => false), (a => 163, b => 167, p => false), (a => 185, b => 189, p => false), (a => 207, b => 211, p => false), (a => 229, b => 233, p => false), (a => 251, b => 255, p => false), (a => 273, b => 277, p => false), (a => 295, b => 299, p => false), (a => 317, b => 321, p => false), (a => 339, b => 343, p => false), (a => 1, b => 5, p => false), (a => 23, b => 27, p => false), (a => 45, b => 49, p => false), (a => 67, b => 71, p => false), (a => 89, b => 93, p => false), (a => 111, b => 115, p => false), (a => 133, b => 137, p => false), (a => 155, b => 159, p => false), (a => 177, b => 181, p => false), (a => 199, b => 203, p => false), (a => 221, b => 225, p => false), (a => 243, b => 247, p => false), (a => 265, b => 269, p => false), (a => 287, b => 291, p => false), (a => 309, b => 313, p => false), (a => 331, b => 335, p => false), (a => 8, b => 12, p => false), (a => 30, b => 34, p => false), (a => 52, b => 56, p => false), (a => 74, b => 78, p => false), (a => 96, b => 100, p => false), (a => 118, b => 122, p => false), (a => 140, b => 144, p => false), (a => 162, b => 166, p => false), (a => 184, b => 188, p => false), (a => 206, b => 210, p => false), (a => 228, b => 232, p => false), (a => 250, b => 254, p => false), (a => 272, b => 276, p => false), (a => 294, b => 298, p => false), (a => 316, b => 320, p => false), (a => 338, b => 342, p => false), (a => 0, b => 4, p => false), (a => 22, b => 26, p => false), (a => 44, b => 48, p => false), (a => 66, b => 70, p => false), (a => 88, b => 92, p => false), (a => 110, b => 114, p => false), (a => 132, b => 136, p => false), (a => 154, b => 158, p => false), (a => 176, b => 180, p => false), (a => 198, b => 202, p => false), (a => 220, b => 224, p => false), (a => 242, b => 246, p => false), (a => 264, b => 268, p => false), (a => 286, b => 290, p => false), (a => 308, b => 312, p => false), (a => 330, b => 334, p => false)),
        ((a    => 4, b => 12, p => false), (a => 26, b => 34, p => false), (a => 48, b => 56, p => false), (a => 70, b => 78, p => false), (a => 92, b => 100, p => false), (a => 114, b => 122, p => false), (a => 136, b => 144, p => false), (a => 158, b => 166, p => false), (a => 180, b => 188, p => false), (a => 202, b => 210, p => false), (a => 224, b => 232, p => false), (a => 246, b => 254, p => false), (a => 268, b => 276, p => false), (a => 290, b => 298, p => false), (a => 312, b => 320, p => false), (a => 334, b => 342, p => false), (a => 17, b => 19, p => false), (a => 39, b => 41, p => false), (a => 61, b => 63, p => false), (a => 83, b => 85, p => false), (a => 105, b => 107, p => false), (a => 127, b => 129, p => false), (a => 149, b => 151, p => false), (a => 171, b => 173, p => false), (a => 193, b => 195, p => false), (a => 215, b => 217, p => false), (a => 237, b => 239, p => false), (a => 259, b => 261, p => false), (a => 281, b => 283, p => false), (a => 303, b => 305, p => false), (a => 325, b => 327, p => false), (a => 347, b => 349, p => false), (a => 6, b => 14, p => false), (a => 28, b => 36, p => false), (a => 50, b => 58, p => false), (a => 72, b => 80, p => false), (a => 94, b => 102, p => false), (a => 116, b => 124, p => false), (a => 138, b => 146, p => false), (a => 160, b => 168, p => false), (a => 182, b => 190, p => false), (a => 204, b => 212, p => false), (a => 226, b => 234, p => false), (a => 248, b => 256, p => false), (a => 270, b => 278, p => false), (a => 292, b => 300, p => false), (a => 314, b => 322, p => false), (a => 336, b => 344, p => false), (a => 2, b => 10, p => false), (a => 24, b => 32, p => false), (a => 46, b => 54, p => false), (a => 68, b => 76, p => false), (a => 90, b => 98, p => false), (a => 112, b => 120, p => false), (a => 134, b => 142, p => false), (a => 156, b => 164, p => false), (a => 178, b => 186, p => false), (a => 200, b => 208, p => false), (a => 222, b => 230, p => false), (a => 244, b => 252, p => false), (a => 266, b => 274, p => false), (a => 288, b => 296, p => false), (a => 310, b => 318, p => false), (a => 332, b => 340, p => false), (a => 11, b => 21, p => false), (a => 33, b => 43, p => false), (a => 55, b => 65, p => false), (a => 77, b => 87, p => false), (a => 99, b => 109, p => false), (a => 121, b => 131, p => false), (a => 143, b => 153, p => false), (a => 165, b => 175, p => false), (a => 187, b => 197, p => false), (a => 209, b => 219, p => false), (a => 231, b => 241, p => false), (a => 253, b => 263, p => false), (a => 275, b => 285, p => false), (a => 297, b => 307, p => false), (a => 319, b => 329, p => false), (a => 341, b => 351, p => false), (a => 5, b => 13, p => false), (a => 27, b => 35, p => false), (a => 49, b => 57, p => false), (a => 71, b => 79, p => false), (a => 93, b => 101, p => false), (a => 115, b => 123, p => false), (a => 137, b => 145, p => false), (a => 159, b => 167, p => false), (a => 181, b => 189, p => false), (a => 203, b => 211, p => false), (a => 225, b => 233, p => false), (a => 247, b => 255, p => false), (a => 269, b => 277, p => false), (a => 291, b => 299, p => false), (a => 313, b => 321, p => false), (a => 335, b => 343, p => false), (a => 9, b => 18, p => false), (a => 31, b => 40, p => false), (a => 53, b => 62, p => false), (a => 75, b => 84, p => false), (a => 97, b => 106, p => false), (a => 119, b => 128, p => false), (a => 141, b => 150, p => false), (a => 163, b => 172, p => false), (a => 185, b => 194, p => false), (a => 207, b => 216, p => false), (a => 229, b => 238, p => false), (a => 251, b => 260, p => false), (a => 273, b => 282, p => false), (a => 295, b => 304, p => false), (a => 317, b => 326, p => false), (a => 339, b => 348, p => false), (a => 0, b => 8, p => false), (a => 22, b => 30, p => false), (a => 44, b => 52, p => false), (a => 66, b => 74, p => false), (a => 88, b => 96, p => false), (a => 110, b => 118, p => false), (a => 132, b => 140, p => false), (a => 154, b => 162, p => false), (a => 176, b => 184, p => false), (a => 198, b => 206, p => false), (a => 220, b => 228, p => false), (a => 242, b => 250, p => false), (a => 264, b => 272, p => false), (a => 286, b => 294, p => false), (a => 308, b => 316, p => false), (a => 330, b => 338, p => false), (a => 3, b => 20, p => false), (a => 25, b => 42, p => false), (a => 47, b => 64, p => false), (a => 69, b => 86, p => false), (a => 91, b => 108, p => false), (a => 113, b => 130, p => false), (a => 135, b => 152, p => false), (a => 157, b => 174, p => false), (a => 179, b => 196, p => false), (a => 201, b => 218, p => false), (a => 223, b => 240, p => false), (a => 245, b => 262, p => false), (a => 267, b => 284, p => false), (a => 289, b => 306, p => false), (a => 311, b => 328, p => false), (a => 333, b => 350, p => false), (a => 1, b => 16, p => false), (a => 23, b => 38, p => false), (a => 45, b => 60, p => false), (a => 67, b => 82, p => false), (a => 89, b => 104, p => false), (a => 111, b => 126, p => false), (a => 133, b => 148, p => false), (a => 155, b => 170, p => false), (a => 177, b => 192, p => false), (a => 199, b => 214, p => false), (a => 221, b => 236, p => false), (a => 243, b => 258, p => false), (a => 265, b => 280, p => false), (a => 287, b => 302, p => false), (a => 309, b => 324, p => false), (a => 331, b => 346, p => false), (a => 7, b => 15, p => false), (a => 29, b => 37, p => false), (a => 51, b => 59, p => false), (a => 73, b => 81, p => false), (a => 95, b => 103, p => false), (a => 117, b => 125, p => false), (a => 139, b => 147, p => false), (a => 161, b => 169, p => false), (a => 183, b => 191, p => false), (a => 205, b => 213, p => false), (a => 227, b => 235, p => false), (a => 249, b => 257, p => false), (a => 271, b => 279, p => false), (a => 293, b => 301, p => false), (a => 315, b => 323, p => false), (a => 337, b => 345, p => false)),
        ((a    => 14, b => 21, p => false), (a => 36, b => 43, p => false), (a => 58, b => 65, p => false), (a => 80, b => 87, p => false), (a => 102, b => 109, p => false), (a => 124, b => 131, p => false), (a => 146, b => 153, p => false), (a => 168, b => 175, p => false), (a => 190, b => 197, p => false), (a => 212, b => 219, p => false), (a => 234, b => 241, p => false), (a => 256, b => 263, p => false), (a => 278, b => 285, p => false), (a => 300, b => 307, p => false), (a => 322, b => 329, p => false), (a => 344, b => 351, p => false), (a => 1, b => 4, p => false), (a => 23, b => 26, p => false), (a => 45, b => 48, p => false), (a => 67, b => 70, p => false), (a => 89, b => 92, p => false), (a => 111, b => 114, p => false), (a => 133, b => 136, p => false), (a => 155, b => 158, p => false), (a => 177, b => 180, p => false), (a => 199, b => 202, p => false), (a => 221, b => 224, p => false), (a => 243, b => 246, p => false), (a => 265, b => 268, p => false), (a => 287, b => 290, p => false), (a => 309, b => 312, p => false), (a => 331, b => 334, p => false), (a => 7, b => 8, p => false), (a => 29, b => 30, p => false), (a => 51, b => 52, p => false), (a => 73, b => 74, p => false), (a => 95, b => 96, p => false), (a => 117, b => 118, p => false), (a => 139, b => 140, p => false), (a => 161, b => 162, p => false), (a => 183, b => 184, p => false), (a => 205, b => 206, p => false), (a => 227, b => 228, p => false), (a => 249, b => 250, p => false), (a => 271, b => 272, p => false), (a => 293, b => 294, p => false), (a => 315, b => 316, p => false), (a => 337, b => 338, p => false), (a => 6, b => 18, p => false), (a => 28, b => 40, p => false), (a => 50, b => 62, p => false), (a => 72, b => 84, p => false), (a => 94, b => 106, p => false), (a => 116, b => 128, p => false), (a => 138, b => 150, p => false), (a => 160, b => 172, p => false), (a => 182, b => 194, p => false), (a => 204, b => 216, p => false), (a => 226, b => 238, p => false), (a => 248, b => 260, p => false), (a => 270, b => 282, p => false), (a => 292, b => 304, p => false), (a => 314, b => 326, p => false), (a => 336, b => 348, p => false), (a => 3, b => 12, p => false), (a => 25, b => 34, p => false), (a => 47, b => 56, p => false), (a => 69, b => 78, p => false), (a => 91, b => 100, p => false), (a => 113, b => 122, p => false), (a => 135, b => 144, p => false), (a => 157, b => 166, p => false), (a => 179, b => 188, p => false), (a => 201, b => 210, p => false), (a => 223, b => 232, p => false), (a => 245, b => 254, p => false), (a => 267, b => 276, p => false), (a => 289, b => 298, p => false), (a => 311, b => 320, p => false), (a => 333, b => 342, p => false), (a => 13, b => 20, p => false), (a => 35, b => 42, p => false), (a => 57, b => 64, p => false), (a => 79, b => 86, p => false), (a => 101, b => 108, p => false), (a => 123, b => 130, p => false), (a => 145, b => 152, p => false), (a => 167, b => 174, p => false), (a => 189, b => 196, p => false), (a => 211, b => 218, p => false), (a => 233, b => 240, p => false), (a => 255, b => 262, p => false), (a => 277, b => 284, p => false), (a => 299, b => 306, p => false), (a => 321, b => 328, p => false), (a => 343, b => 350, p => false), (a => 10, b => 19, p => false), (a => 32, b => 41, p => false), (a => 54, b => 63, p => false), (a => 76, b => 85, p => false), (a => 98, b => 107, p => false), (a => 120, b => 129, p => false), (a => 142, b => 151, p => false), (a => 164, b => 173, p => false), (a => 186, b => 195, p => false), (a => 208, b => 217, p => false), (a => 230, b => 239, p => false), (a => 252, b => 261, p => false), (a => 274, b => 283, p => false), (a => 296, b => 305, p => false), (a => 318, b => 327, p => false), (a => 340, b => 349, p => false), (a => 2, b => 9, p => false), (a => 24, b => 31, p => false), (a => 46, b => 53, p => false), (a => 68, b => 75, p => false), (a => 90, b => 97, p => false), (a => 112, b => 119, p => false), (a => 134, b => 141, p => false), (a => 156, b => 163, p => false), (a => 178, b => 185, p => false), (a => 200, b => 207, p => false), (a => 222, b => 229, p => false), (a => 244, b => 251, p => false), (a => 266, b => 273, p => false), (a => 288, b => 295, p => false), (a => 310, b => 317, p => false), (a => 332, b => 339, p => false), (a => 5, b => 17, p => false), (a => 27, b => 39, p => false), (a => 49, b => 61, p => false), (a => 71, b => 83, p => false), (a => 93, b => 105, p => false), (a => 115, b => 127, p => false), (a => 137, b => 149, p => false), (a => 159, b => 171, p => false), (a => 181, b => 193, p => false), (a => 203, b => 215, p => false), (a => 225, b => 237, p => false), (a => 247, b => 259, p => false), (a => 269, b => 281, p => false), (a => 291, b => 303, p => false), (a => 313, b => 325, p => false), (a => 335, b => 347, p => false), (a => 11, b => 16, p => false), (a => 33, b => 38, p => false), (a => 55, b => 60, p => false), (a => 77, b => 82, p => false), (a => 99, b => 104, p => false), (a => 121, b => 126, p => false), (a => 143, b => 148, p => false), (a => 165, b => 170, p => false), (a => 187, b => 192, p => false), (a => 209, b => 214, p => false), (a => 231, b => 236, p => false), (a => 253, b => 258, p => false), (a => 275, b => 280, p => false), (a => 297, b => 302, p => false), (a => 319, b => 324, p => false), (a => 341, b => 346, p => false), (a => 0, b => 345, p => true), (a => 15, b => 330, p => true), (a => 22, b => 323, p => true), (a => 37, b => 308, p => true), (a => 44, b => 301, p => true), (a => 59, b => 286, p => true), (a => 66, b => 279, p => true), (a => 81, b => 264, p => true), (a => 88, b => 257, p => true), (a => 103, b => 242, p => true), (a => 110, b => 235, p => true), (a => 125, b => 220, p => true), (a => 132, b => 213, p => true), (a => 147, b => 198, p => true), (a => 154, b => 191, p => true), (a => 169, b => 176, p => true)),
        ((a    => 0, b => 1, p => false), (a => 22, b => 23, p => false), (a => 44, b => 45, p => false), (a => 66, b => 67, p => false), (a => 88, b => 89, p => false), (a => 110, b => 111, p => false), (a => 132, b => 133, p => false), (a => 154, b => 155, p => false), (a => 176, b => 177, p => false), (a => 198, b => 199, p => false), (a => 220, b => 221, p => false), (a => 242, b => 243, p => false), (a => 264, b => 265, p => false), (a => 286, b => 287, p => false), (a => 308, b => 309, p => false), (a => 330, b => 331, p => false), (a => 15, b => 21, p => false), (a => 37, b => 43, p => false), (a => 59, b => 65, p => false), (a => 81, b => 87, p => false), (a => 103, b => 109, p => false), (a => 125, b => 131, p => false), (a => 147, b => 153, p => false), (a => 169, b => 175, p => false), (a => 191, b => 197, p => false), (a => 213, b => 219, p => false), (a => 235, b => 241, p => false), (a => 257, b => 263, p => false), (a => 279, b => 285, p => false), (a => 301, b => 307, p => false), (a => 323, b => 329, p => false), (a => 345, b => 351, p => false), (a => 3, b => 9, p => false), (a => 25, b => 31, p => false), (a => 47, b => 53, p => false), (a => 69, b => 75, p => false), (a => 91, b => 97, p => false), (a => 113, b => 119, p => false), (a => 135, b => 141, p => false), (a => 157, b => 163, p => false), (a => 179, b => 185, p => false), (a => 201, b => 207, p => false), (a => 223, b => 229, p => false), (a => 245, b => 251, p => false), (a => 267, b => 273, p => false), (a => 289, b => 295, p => false), (a => 311, b => 317, p => false), (a => 333, b => 339, p => false), (a => 13, b => 18, p => false), (a => 35, b => 40, p => false), (a => 57, b => 62, p => false), (a => 79, b => 84, p => false), (a => 101, b => 106, p => false), (a => 123, b => 128, p => false), (a => 145, b => 150, p => false), (a => 167, b => 172, p => false), (a => 189, b => 194, p => false), (a => 211, b => 216, p => false), (a => 233, b => 238, p => false), (a => 255, b => 260, p => false), (a => 277, b => 282, p => false), (a => 299, b => 304, p => false), (a => 321, b => 326, p => false), (a => 343, b => 348, p => false), (a => 5, b => 7, p => false), (a => 27, b => 29, p => false), (a => 49, b => 51, p => false), (a => 71, b => 73, p => false), (a => 93, b => 95, p => false), (a => 115, b => 117, p => false), (a => 137, b => 139, p => false), (a => 159, b => 161, p => false), (a => 181, b => 183, p => false), (a => 203, b => 205, p => false), (a => 225, b => 227, p => false), (a => 247, b => 249, p => false), (a => 269, b => 271, p => false), (a => 291, b => 293, p => false), (a => 313, b => 315, p => false), (a => 335, b => 337, p => false), (a => 8, b => 19, p => false), (a => 30, b => 41, p => false), (a => 52, b => 63, p => false), (a => 74, b => 85, p => false), (a => 96, b => 107, p => false), (a => 118, b => 129, p => false), (a => 140, b => 151, p => false), (a => 162, b => 173, p => false), (a => 184, b => 195, p => false), (a => 206, b => 217, p => false), (a => 228, b => 239, p => false), (a => 250, b => 261, p => false), (a => 272, b => 283, p => false), (a => 294, b => 305, p => false), (a => 316, b => 327, p => false), (a => 338, b => 349, p => false), (a => 12, b => 16, p => false), (a => 34, b => 38, p => false), (a => 56, b => 60, p => false), (a => 78, b => 82, p => false), (a => 100, b => 104, p => false), (a => 122, b => 126, p => false), (a => 144, b => 148, p => false), (a => 166, b => 170, p => false), (a => 188, b => 192, p => false), (a => 210, b => 214, p => false), (a => 232, b => 236, p => false), (a => 254, b => 258, p => false), (a => 276, b => 280, p => false), (a => 298, b => 302, p => false), (a => 320, b => 324, p => false), (a => 342, b => 346, p => false), (a => 6, b => 11, p => false), (a => 28, b => 33, p => false), (a => 50, b => 55, p => false), (a => 72, b => 77, p => false), (a => 94, b => 99, p => false), (a => 116, b => 121, p => false), (a => 138, b => 143, p => false), (a => 160, b => 165, p => false), (a => 182, b => 187, p => false), (a => 204, b => 209, p => false), (a => 226, b => 231, p => false), (a => 248, b => 253, p => false), (a => 270, b => 275, p => false), (a => 292, b => 297, p => false), (a => 314, b => 319, p => false), (a => 336, b => 341, p => false), (a => 14, b => 17, p => false), (a => 36, b => 39, p => false), (a => 58, b => 61, p => false), (a => 80, b => 83, p => false), (a => 102, b => 105, p => false), (a => 124, b => 127, p => false), (a => 146, b => 149, p => false), (a => 168, b => 171, p => false), (a => 190, b => 193, p => false), (a => 212, b => 215, p => false), (a => 234, b => 237, p => false), (a => 256, b => 259, p => false), (a => 278, b => 281, p => false), (a => 300, b => 303, p => false), (a => 322, b => 325, p => false), (a => 344, b => 347, p => false), (a => 4, b => 10, p => false), (a => 26, b => 32, p => false), (a => 48, b => 54, p => false), (a => 70, b => 76, p => false), (a => 92, b => 98, p => false), (a => 114, b => 120, p => false), (a => 136, b => 142, p => false), (a => 158, b => 164, p => false), (a => 180, b => 186, p => false), (a => 202, b => 208, p => false), (a => 224, b => 230, p => false), (a => 246, b => 252, p => false), (a => 268, b => 274, p => false), (a => 290, b => 296, p => false), (a => 312, b => 318, p => false), (a => 334, b => 340, p => false), (a => 2, b => 350, p => true), (a => 20, b => 332, p => true), (a => 24, b => 328, p => true), (a => 42, b => 310, p => true), (a => 46, b => 306, p => true), (a => 64, b => 288, p => true), (a => 68, b => 284, p => true), (a => 86, b => 266, p => true), (a => 90, b => 262, p => true), (a => 108, b => 244, p => true), (a => 112, b => 240, p => true), (a => 130, b => 222, p => true), (a => 134, b => 218, p => true), (a => 152, b => 200, p => true), (a => 156, b => 196, p => true), (a => 174, b => 178, p => true)),
        ((a    => 1, b => 5, p => false), (a => 23, b => 27, p => false), (a => 45, b => 49, p => false), (a => 67, b => 71, p => false), (a => 89, b => 93, p => false), (a => 111, b => 115, p => false), (a => 133, b => 137, p => false), (a => 155, b => 159, p => false), (a => 177, b => 181, p => false), (a => 199, b => 203, p => false), (a => 221, b => 225, p => false), (a => 243, b => 247, p => false), (a => 265, b => 269, p => false), (a => 287, b => 291, p => false), (a => 309, b => 313, p => false), (a => 331, b => 335, p => false), (a => 7, b => 9, p => false), (a => 29, b => 31, p => false), (a => 51, b => 53, p => false), (a => 73, b => 75, p => false), (a => 95, b => 97, p => false), (a => 117, b => 119, p => false), (a => 139, b => 141, p => false), (a => 161, b => 163, p => false), (a => 183, b => 185, p => false), (a => 205, b => 207, p => false), (a => 227, b => 229, p => false), (a => 249, b => 251, p => false), (a => 271, b => 273, p => false), (a => 293, b => 295, p => false), (a => 315, b => 317, p => false), (a => 337, b => 339, p => false), (a => 10, b => 11, p => false), (a => 32, b => 33, p => false), (a => 54, b => 55, p => false), (a => 76, b => 77, p => false), (a => 98, b => 99, p => false), (a => 120, b => 121, p => false), (a => 142, b => 143, p => false), (a => 164, b => 165, p => false), (a => 186, b => 187, p => false), (a => 208, b => 209, p => false), (a => 230, b => 231, p => false), (a => 252, b => 253, p => false), (a => 274, b => 275, p => false), (a => 296, b => 297, p => false), (a => 318, b => 319, p => false), (a => 340, b => 341, p => false), (a => 12, b => 14, p => false), (a => 34, b => 36, p => false), (a => 56, b => 58, p => false), (a => 78, b => 80, p => false), (a => 100, b => 102, p => false), (a => 122, b => 124, p => false), (a => 144, b => 146, p => false), (a => 166, b => 168, p => false), (a => 188, b => 190, p => false), (a => 210, b => 212, p => false), (a => 232, b => 234, p => false), (a => 254, b => 256, p => false), (a => 276, b => 278, p => false), (a => 298, b => 300, p => false), (a => 320, b => 322, p => false), (a => 342, b => 344, p => false), (a => 16, b => 17, p => false), (a => 38, b => 39, p => false), (a => 60, b => 61, p => false), (a => 82, b => 83, p => false), (a => 104, b => 105, p => false), (a => 126, b => 127, p => false), (a => 148, b => 149, p => false), (a => 170, b => 171, p => false), (a => 192, b => 193, p => false), (a => 214, b => 215, p => false), (a => 236, b => 237, p => false), (a => 258, b => 259, p => false), (a => 280, b => 281, p => false), (a => 302, b => 303, p => false), (a => 324, b => 325, p => false), (a => 346, b => 347, p => false), (a => 18, b => 20, p => false), (a => 40, b => 42, p => false), (a => 62, b => 64, p => false), (a => 84, b => 86, p => false), (a => 106, b => 108, p => false), (a => 128, b => 130, p => false), (a => 150, b => 152, p => false), (a => 172, b => 174, p => false), (a => 194, b => 196, p => false), (a => 216, b => 218, p => false), (a => 238, b => 240, p => false), (a => 260, b => 262, p => false), (a => 282, b => 284, p => false), (a => 304, b => 306, p => false), (a => 326, b => 328, p => false), (a => 348, b => 350, p => false), (a => 2, b => 3, p => false), (a => 24, b => 25, p => false), (a => 46, b => 47, p => false), (a => 68, b => 69, p => false), (a => 90, b => 91, p => false), (a => 112, b => 113, p => false), (a => 134, b => 135, p => false), (a => 156, b => 157, p => false), (a => 178, b => 179, p => false), (a => 200, b => 201, p => false), (a => 222, b => 223, p => false), (a => 244, b => 245, p => false), (a => 266, b => 267, p => false), (a => 288, b => 289, p => false), (a => 310, b => 311, p => false), (a => 332, b => 333, p => false), (a => 4, b => 6, p => false), (a => 26, b => 28, p => false), (a => 48, b => 50, p => false), (a => 70, b => 72, p => false), (a => 92, b => 94, p => false), (a => 114, b => 116, p => false), (a => 136, b => 138, p => false), (a => 158, b => 160, p => false), (a => 180, b => 182, p => false), (a => 202, b => 204, p => false), (a => 224, b => 226, p => false), (a => 246, b => 248, p => false), (a => 268, b => 270, p => false), (a => 290, b => 292, p => false), (a => 312, b => 314, p => false), (a => 334, b => 336, p => false), (a => 8, b => 13, p => false), (a => 30, b => 35, p => false), (a => 52, b => 57, p => false), (a => 74, b => 79, p => false), (a => 96, b => 101, p => false), (a => 118, b => 123, p => false), (a => 140, b => 145, p => false), (a => 162, b => 167, p => false), (a => 184, b => 189, p => false), (a => 206, b => 211, p => false), (a => 228, b => 233, p => false), (a => 250, b => 255, p => false), (a => 272, b => 277, p => false), (a => 294, b => 299, p => false), (a => 316, b => 321, p => false), (a => 338, b => 343, p => false), (a => 15, b => 19, p => false), (a => 37, b => 41, p => false), (a => 59, b => 63, p => false), (a => 81, b => 85, p => false), (a => 103, b => 107, p => false), (a => 125, b => 129, p => false), (a => 147, b => 151, p => false), (a => 169, b => 173, p => false), (a => 191, b => 195, p => false), (a => 213, b => 217, p => false), (a => 235, b => 239, p => false), (a => 257, b => 261, p => false), (a => 279, b => 283, p => false), (a => 301, b => 305, p => false), (a => 323, b => 327, p => false), (a => 345, b => 349, p => false), (a => 0, b => 22, p => false), (a => 44, b => 66, p => false), (a => 88, b => 110, p => false), (a => 132, b => 154, p => false), (a => 176, b => 198, p => false), (a => 220, b => 242, p => false), (a => 264, b => 286, p => false), (a => 308, b => 330, p => false), (a => 21, b => 351, p => true), (a => 43, b => 329, p => true), (a => 65, b => 307, p => true), (a => 87, b => 285, p => true), (a => 109, b => 263, p => true), (a => 131, b => 241, p => true), (a => 153, b => 219, p => true), (a => 175, b => 197, p => true)),
        ((a    => 1, b => 2, p => false), (a => 23, b => 24, p => false), (a => 45, b => 46, p => false), (a => 67, b => 68, p => false), (a => 89, b => 90, p => false), (a => 111, b => 112, p => false), (a => 133, b => 134, p => false), (a => 155, b => 156, p => false), (a => 177, b => 178, p => false), (a => 199, b => 200, p => false), (a => 221, b => 222, p => false), (a => 243, b => 244, p => false), (a => 265, b => 266, p => false), (a => 287, b => 288, p => false), (a => 309, b => 310, p => false), (a => 331, b => 332, p => false), (a => 4, b => 5, p => false), (a => 26, b => 27, p => false), (a => 48, b => 49, p => false), (a => 70, b => 71, p => false), (a => 92, b => 93, p => false), (a => 114, b => 115, p => false), (a => 136, b => 137, p => false), (a => 158, b => 159, p => false), (a => 180, b => 181, p => false), (a => 202, b => 203, p => false), (a => 224, b => 225, p => false), (a => 246, b => 247, p => false), (a => 268, b => 269, p => false), (a => 290, b => 291, p => false), (a => 312, b => 313, p => false), (a => 334, b => 335, p => false), (a => 7, b => 10, p => false), (a => 29, b => 32, p => false), (a => 51, b => 54, p => false), (a => 73, b => 76, p => false), (a => 95, b => 98, p => false), (a => 117, b => 120, p => false), (a => 139, b => 142, p => false), (a => 161, b => 164, p => false), (a => 183, b => 186, p => false), (a => 205, b => 208, p => false), (a => 227, b => 230, p => false), (a => 249, b => 252, p => false), (a => 271, b => 274, p => false), (a => 293, b => 296, p => false), (a => 315, b => 318, p => false), (a => 337, b => 340, p => false), (a => 13, b => 14, p => false), (a => 35, b => 36, p => false), (a => 57, b => 58, p => false), (a => 79, b => 80, p => false), (a => 101, b => 102, p => false), (a => 123, b => 124, p => false), (a => 145, b => 146, p => false), (a => 167, b => 168, p => false), (a => 189, b => 190, p => false), (a => 211, b => 212, p => false), (a => 233, b => 234, p => false), (a => 255, b => 256, p => false), (a => 277, b => 278, p => false), (a => 299, b => 300, p => false), (a => 321, b => 322, p => false), (a => 343, b => 344, p => false), (a => 16, b => 18, p => false), (a => 38, b => 40, p => false), (a => 60, b => 62, p => false), (a => 82, b => 84, p => false), (a => 104, b => 106, p => false), (a => 126, b => 128, p => false), (a => 148, b => 150, p => false), (a => 170, b => 172, p => false), (a => 192, b => 194, p => false), (a => 214, b => 216, p => false), (a => 236, b => 238, p => false), (a => 258, b => 260, p => false), (a => 280, b => 282, p => false), (a => 302, b => 304, p => false), (a => 324, b => 326, p => false), (a => 346, b => 348, p => false), (a => 19, b => 20, p => false), (a => 41, b => 42, p => false), (a => 63, b => 64, p => false), (a => 85, b => 86, p => false), (a => 107, b => 108, p => false), (a => 129, b => 130, p => false), (a => 151, b => 152, p => false), (a => 173, b => 174, p => false), (a => 195, b => 196, p => false), (a => 217, b => 218, p => false), (a => 239, b => 240, p => false), (a => 261, b => 262, p => false), (a => 283, b => 284, p => false), (a => 305, b => 306, p => false), (a => 327, b => 328, p => false), (a => 349, b => 350, p => false), (a => 3, b => 6, p => false), (a => 25, b => 28, p => false), (a => 47, b => 50, p => false), (a => 69, b => 72, p => false), (a => 91, b => 94, p => false), (a => 113, b => 116, p => false), (a => 135, b => 138, p => false), (a => 157, b => 160, p => false), (a => 179, b => 182, p => false), (a => 201, b => 204, p => false), (a => 223, b => 226, p => false), (a => 245, b => 248, p => false), (a => 267, b => 270, p => false), (a => 289, b => 292, p => false), (a => 311, b => 314, p => false), (a => 333, b => 336, p => false), (a => 8, b => 12, p => false), (a => 30, b => 34, p => false), (a => 52, b => 56, p => false), (a => 74, b => 78, p => false), (a => 96, b => 100, p => false), (a => 118, b => 122, p => false), (a => 140, b => 144, p => false), (a => 162, b => 166, p => false), (a => 184, b => 188, p => false), (a => 206, b => 210, p => false), (a => 228, b => 232, p => false), (a => 250, b => 254, p => false), (a => 272, b => 276, p => false), (a => 294, b => 298, p => false), (a => 316, b => 320, p => false), (a => 338, b => 342, p => false), (a => 15, b => 17, p => false), (a => 37, b => 39, p => false), (a => 59, b => 61, p => false), (a => 81, b => 83, p => false), (a => 103, b => 105, p => false), (a => 125, b => 127, p => false), (a => 147, b => 149, p => false), (a => 169, b => 171, p => false), (a => 191, b => 193, p => false), (a => 213, b => 215, p => false), (a => 235, b => 237, p => false), (a => 257, b => 259, p => false), (a => 279, b => 281, p => false), (a => 301, b => 303, p => false), (a => 323, b => 325, p => false), (a => 345, b => 347, p => false), (a => 9, b => 11, p => false), (a => 31, b => 33, p => false), (a => 53, b => 55, p => false), (a => 75, b => 77, p => false), (a => 97, b => 99, p => false), (a => 119, b => 121, p => false), (a => 141, b => 143, p => false), (a => 163, b => 165, p => false), (a => 185, b => 187, p => false), (a => 207, b => 209, p => false), (a => 229, b => 231, p => false), (a => 251, b => 253, p => false), (a => 273, b => 275, p => false), (a => 295, b => 297, p => false), (a => 317, b => 319, p => false), (a => 339, b => 341, p => false), (a => 0, b => 44, p => false), (a => 88, b => 132, p => false), (a => 176, b => 220, p => false), (a => 264, b => 308, p => false), (a => 21, b => 351, p => true), (a => 22, b => 330, p => true), (a => 43, b => 329, p => true), (a => 65, b => 307, p => true), (a => 66, b => 286, p => true), (a => 87, b => 285, p => true), (a => 109, b => 263, p => true), (a => 110, b => 242, p => true), (a => 131, b => 241, p => true), (a => 153, b => 219, p => true), (a => 154, b => 198, p => true), (a => 175, b => 197, p => true)),
        ((a    => 2, b => 3, p => false), (a => 24, b => 25, p => false), (a => 46, b => 47, p => false), (a => 68, b => 69, p => false), (a => 90, b => 91, p => false), (a => 112, b => 113, p => false), (a => 134, b => 135, p => false), (a => 156, b => 157, p => false), (a => 178, b => 179, p => false), (a => 200, b => 201, p => false), (a => 222, b => 223, p => false), (a => 244, b => 245, p => false), (a => 266, b => 267, p => false), (a => 288, b => 289, p => false), (a => 310, b => 311, p => false), (a => 332, b => 333, p => false), (a => 5, b => 7, p => false), (a => 27, b => 29, p => false), (a => 49, b => 51, p => false), (a => 71, b => 73, p => false), (a => 93, b => 95, p => false), (a => 115, b => 117, p => false), (a => 137, b => 139, p => false), (a => 159, b => 161, p => false), (a => 181, b => 183, p => false), (a => 203, b => 205, p => false), (a => 225, b => 227, p => false), (a => 247, b => 249, p => false), (a => 269, b => 271, p => false), (a => 291, b => 293, p => false), (a => 313, b => 315, p => false), (a => 335, b => 337, p => false), (a => 9, b => 10, p => false), (a => 31, b => 32, p => false), (a => 53, b => 54, p => false), (a => 75, b => 76, p => false), (a => 97, b => 98, p => false), (a => 119, b => 120, p => false), (a => 141, b => 142, p => false), (a => 163, b => 164, p => false), (a => 185, b => 186, p => false), (a => 207, b => 208, p => false), (a => 229, b => 230, p => false), (a => 251, b => 252, p => false), (a => 273, b => 274, p => false), (a => 295, b => 296, p => false), (a => 317, b => 318, p => false), (a => 339, b => 340, p => false), (a => 12, b => 13, p => false), (a => 34, b => 35, p => false), (a => 56, b => 57, p => false), (a => 78, b => 79, p => false), (a => 100, b => 101, p => false), (a => 122, b => 123, p => false), (a => 144, b => 145, p => false), (a => 166, b => 167, p => false), (a => 188, b => 189, p => false), (a => 210, b => 211, p => false), (a => 232, b => 233, p => false), (a => 254, b => 255, p => false), (a => 276, b => 277, p => false), (a => 298, b => 299, p => false), (a => 320, b => 321, p => false), (a => 342, b => 343, p => false), (a => 14, b => 15, p => false), (a => 36, b => 37, p => false), (a => 58, b => 59, p => false), (a => 80, b => 81, p => false), (a => 102, b => 103, p => false), (a => 124, b => 125, p => false), (a => 146, b => 147, p => false), (a => 168, b => 169, p => false), (a => 190, b => 191, p => false), (a => 212, b => 213, p => false), (a => 234, b => 235, p => false), (a => 256, b => 257, p => false), (a => 278, b => 279, p => false), (a => 300, b => 301, p => false), (a => 322, b => 323, p => false), (a => 344, b => 345, p => false), (a => 18, b => 19, p => false), (a => 40, b => 41, p => false), (a => 62, b => 63, p => false), (a => 84, b => 85, p => false), (a => 106, b => 107, p => false), (a => 128, b => 129, p => false), (a => 150, b => 151, p => false), (a => 172, b => 173, p => false), (a => 194, b => 195, p => false), (a => 216, b => 217, p => false), (a => 238, b => 239, p => false), (a => 260, b => 261, p => false), (a => 282, b => 283, p => false), (a => 304, b => 305, p => false), (a => 326, b => 327, p => false), (a => 348, b => 349, p => false), (a => 6, b => 8, p => false), (a => 28, b => 30, p => false), (a => 50, b => 52, p => false), (a => 72, b => 74, p => false), (a => 94, b => 96, p => false), (a => 116, b => 118, p => false), (a => 138, b => 140, p => false), (a => 160, b => 162, p => false), (a => 182, b => 184, p => false), (a => 204, b => 206, p => false), (a => 226, b => 228, p => false), (a => 248, b => 250, p => false), (a => 270, b => 272, p => false), (a => 292, b => 294, p => false), (a => 314, b => 316, p => false), (a => 336, b => 338, p => false), (a => 11, b => 16, p => false), (a => 33, b => 38, p => false), (a => 55, b => 60, p => false), (a => 77, b => 82, p => false), (a => 99, b => 104, p => false), (a => 121, b => 126, p => false), (a => 143, b => 148, p => false), (a => 165, b => 170, p => false), (a => 187, b => 192, p => false), (a => 209, b => 214, p => false), (a => 231, b => 236, p => false), (a => 253, b => 258, p => false), (a => 275, b => 280, p => false), (a => 297, b => 302, p => false), (a => 319, b => 324, p => false), (a => 341, b => 346, p => false), (a => 1, b => 23, p => false), (a => 45, b => 67, p => false), (a => 89, b => 111, p => false), (a => 133, b => 155, p => false), (a => 177, b => 199, p => false), (a => 221, b => 243, p => false), (a => 265, b => 287, p => false), (a => 309, b => 331, p => false), (a => 0, b => 88, p => false), (a => 176, b => 264, p => false), (a => 4, b => 351, p => true), (a => 17, b => 350, p => true), (a => 20, b => 347, p => true), (a => 21, b => 334, p => true), (a => 22, b => 330, p => true), (a => 26, b => 329, p => true), (a => 39, b => 328, p => true), (a => 42, b => 325, p => true), (a => 43, b => 312, p => true), (a => 44, b => 308, p => true), (a => 48, b => 307, p => true), (a => 61, b => 306, p => true), (a => 64, b => 303, p => true), (a => 65, b => 290, p => true), (a => 66, b => 286, p => true), (a => 70, b => 285, p => true), (a => 83, b => 284, p => true), (a => 86, b => 281, p => true), (a => 87, b => 268, p => true), (a => 92, b => 263, p => true), (a => 105, b => 262, p => true), (a => 108, b => 259, p => true), (a => 109, b => 246, p => true), (a => 110, b => 242, p => true), (a => 114, b => 241, p => true), (a => 127, b => 240, p => true), (a => 130, b => 237, p => true), (a => 131, b => 224, p => true), (a => 132, b => 220, p => true), (a => 136, b => 219, p => true), (a => 149, b => 218, p => true), (a => 152, b => 215, p => true), (a => 153, b => 202, p => true), (a => 154, b => 198, p => true), (a => 158, b => 197, p => true), (a => 171, b => 196, p => true), (a => 174, b => 193, p => true), (a => 175, b => 180, p => true)),
        ((a    => 2, b => 4, p => false), (a => 24, b => 26, p => false), (a => 46, b => 48, p => false), (a => 68, b => 70, p => false), (a => 90, b => 92, p => false), (a => 112, b => 114, p => false), (a => 134, b => 136, p => false), (a => 156, b => 158, p => false), (a => 178, b => 180, p => false), (a => 200, b => 202, p => false), (a => 222, b => 224, p => false), (a => 244, b => 246, p => false), (a => 266, b => 268, p => false), (a => 288, b => 290, p => false), (a => 310, b => 312, p => false), (a => 332, b => 334, p => false), (a => 6, b => 7, p => false), (a => 28, b => 29, p => false), (a => 50, b => 51, p => false), (a => 72, b => 73, p => false), (a => 94, b => 95, p => false), (a => 116, b => 117, p => false), (a => 138, b => 139, p => false), (a => 160, b => 161, p => false), (a => 182, b => 183, p => false), (a => 204, b => 205, p => false), (a => 226, b => 227, p => false), (a => 248, b => 249, p => false), (a => 270, b => 271, p => false), (a => 292, b => 293, p => false), (a => 314, b => 315, p => false), (a => 336, b => 337, p => false), (a => 8, b => 9, p => false), (a => 30, b => 31, p => false), (a => 52, b => 53, p => false), (a => 74, b => 75, p => false), (a => 96, b => 97, p => false), (a => 118, b => 119, p => false), (a => 140, b => 141, p => false), (a => 162, b => 163, p => false), (a => 184, b => 185, p => false), (a => 206, b => 207, p => false), (a => 228, b => 229, p => false), (a => 250, b => 251, p => false), (a => 272, b => 273, p => false), (a => 294, b => 295, p => false), (a => 316, b => 317, p => false), (a => 338, b => 339, p => false), (a => 10, b => 12, p => false), (a => 32, b => 34, p => false), (a => 54, b => 56, p => false), (a => 76, b => 78, p => false), (a => 98, b => 100, p => false), (a => 120, b => 122, p => false), (a => 142, b => 144, p => false), (a => 164, b => 166, p => false), (a => 186, b => 188, p => false), (a => 208, b => 210, p => false), (a => 230, b => 232, p => false), (a => 252, b => 254, p => false), (a => 274, b => 276, p => false), (a => 296, b => 298, p => false), (a => 318, b => 320, p => false), (a => 340, b => 342, p => false), (a => 14, b => 16, p => false), (a => 36, b => 38, p => false), (a => 58, b => 60, p => false), (a => 80, b => 82, p => false), (a => 102, b => 104, p => false), (a => 124, b => 126, p => false), (a => 146, b => 148, p => false), (a => 168, b => 170, p => false), (a => 190, b => 192, p => false), (a => 212, b => 214, p => false), (a => 234, b => 236, p => false), (a => 256, b => 258, p => false), (a => 278, b => 280, p => false), (a => 300, b => 302, p => false), (a => 322, b => 324, p => false), (a => 344, b => 346, p => false), (a => 3, b => 5, p => false), (a => 25, b => 27, p => false), (a => 47, b => 49, p => false), (a => 69, b => 71, p => false), (a => 91, b => 93, p => false), (a => 113, b => 115, p => false), (a => 135, b => 137, p => false), (a => 157, b => 159, p => false), (a => 179, b => 181, p => false), (a => 201, b => 203, p => false), (a => 223, b => 225, p => false), (a => 245, b => 247, p => false), (a => 267, b => 269, p => false), (a => 289, b => 291, p => false), (a => 311, b => 313, p => false), (a => 333, b => 335, p => false), (a => 11, b => 13, p => false), (a => 33, b => 35, p => false), (a => 55, b => 57, p => false), (a => 77, b => 79, p => false), (a => 99, b => 101, p => false), (a => 121, b => 123, p => false), (a => 143, b => 145, p => false), (a => 165, b => 167, p => false), (a => 187, b => 189, p => false), (a => 209, b => 211, p => false), (a => 231, b => 233, p => false), (a => 253, b => 255, p => false), (a => 275, b => 277, p => false), (a => 297, b => 299, p => false), (a => 319, b => 321, p => false), (a => 341, b => 343, p => false), (a => 15, b => 18, p => false), (a => 37, b => 40, p => false), (a => 59, b => 62, p => false), (a => 81, b => 84, p => false), (a => 103, b => 106, p => false), (a => 125, b => 128, p => false), (a => 147, b => 150, p => false), (a => 169, b => 172, p => false), (a => 191, b => 194, p => false), (a => 213, b => 216, p => false), (a => 235, b => 238, p => false), (a => 257, b => 260, p => false), (a => 279, b => 282, p => false), (a => 301, b => 304, p => false), (a => 323, b => 326, p => false), (a => 345, b => 348, p => false), (a => 0, b => 176, p => false), (a => 1, b => 351, p => true), (a => 17, b => 350, p => true), (a => 19, b => 349, p => true), (a => 20, b => 347, p => true), (a => 21, b => 331, p => true), (a => 22, b => 330, p => true), (a => 23, b => 329, p => true), (a => 39, b => 328, p => true), (a => 41, b => 327, p => true), (a => 42, b => 325, p => true), (a => 43, b => 309, p => true), (a => 44, b => 308, p => true), (a => 45, b => 307, p => true), (a => 61, b => 306, p => true), (a => 63, b => 305, p => true), (a => 64, b => 303, p => true), (a => 65, b => 287, p => true), (a => 66, b => 286, p => true), (a => 67, b => 285, p => true), (a => 83, b => 284, p => true), (a => 85, b => 283, p => true), (a => 86, b => 281, p => true), (a => 87, b => 265, p => true), (a => 88, b => 264, p => true), (a => 89, b => 263, p => true), (a => 105, b => 262, p => true), (a => 107, b => 261, p => true), (a => 108, b => 259, p => true), (a => 109, b => 243, p => true), (a => 110, b => 242, p => true), (a => 111, b => 241, p => true), (a => 127, b => 240, p => true), (a => 129, b => 239, p => true), (a => 130, b => 237, p => true), (a => 131, b => 221, p => true), (a => 132, b => 220, p => true), (a => 133, b => 219, p => true), (a => 149, b => 218, p => true), (a => 151, b => 217, p => true), (a => 152, b => 215, p => true), (a => 153, b => 199, p => true), (a => 154, b => 198, p => true), (a => 155, b => 197, p => true), (a => 171, b => 196, p => true), (a => 173, b => 195, p => true), (a => 174, b => 193, p => true), (a => 175, b => 177, p => true)),
        ((a    => 3, b => 4, p => false), (a => 25, b => 26, p => false), (a => 47, b => 48, p => false), (a => 69, b => 70, p => false), (a => 91, b => 92, p => false), (a => 113, b => 114, p => false), (a => 135, b => 136, p => false), (a => 157, b => 158, p => false), (a => 179, b => 180, p => false), (a => 201, b => 202, p => false), (a => 223, b => 224, p => false), (a => 245, b => 246, p => false), (a => 267, b => 268, p => false), (a => 289, b => 290, p => false), (a => 311, b => 312, p => false), (a => 333, b => 334, p => false), (a => 5, b => 6, p => false), (a => 27, b => 28, p => false), (a => 49, b => 50, p => false), (a => 71, b => 72, p => false), (a => 93, b => 94, p => false), (a => 115, b => 116, p => false), (a => 137, b => 138, p => false), (a => 159, b => 160, p => false), (a => 181, b => 182, p => false), (a => 203, b => 204, p => false), (a => 225, b => 226, p => false), (a => 247, b => 248, p => false), (a => 269, b => 270, p => false), (a => 291, b => 292, p => false), (a => 313, b => 314, p => false), (a => 335, b => 336, p => false), (a => 7, b => 8, p => false), (a => 29, b => 30, p => false), (a => 51, b => 52, p => false), (a => 73, b => 74, p => false), (a => 95, b => 96, p => false), (a => 117, b => 118, p => false), (a => 139, b => 140, p => false), (a => 161, b => 162, p => false), (a => 183, b => 184, p => false), (a => 205, b => 206, p => false), (a => 227, b => 228, p => false), (a => 249, b => 250, p => false), (a => 271, b => 272, p => false), (a => 293, b => 294, p => false), (a => 315, b => 316, p => false), (a => 337, b => 338, p => false), (a => 9, b => 10, p => false), (a => 31, b => 32, p => false), (a => 53, b => 54, p => false), (a => 75, b => 76, p => false), (a => 97, b => 98, p => false), (a => 119, b => 120, p => false), (a => 141, b => 142, p => false), (a => 163, b => 164, p => false), (a => 185, b => 186, p => false), (a => 207, b => 208, p => false), (a => 229, b => 230, p => false), (a => 251, b => 252, p => false), (a => 273, b => 274, p => false), (a => 295, b => 296, p => false), (a => 317, b => 318, p => false), (a => 339, b => 340, p => false), (a => 11, b => 12, p => false), (a => 33, b => 34, p => false), (a => 55, b => 56, p => false), (a => 77, b => 78, p => false), (a => 99, b => 100, p => false), (a => 121, b => 122, p => false), (a => 143, b => 144, p => false), (a => 165, b => 166, p => false), (a => 187, b => 188, p => false), (a => 209, b => 210, p => false), (a => 231, b => 232, p => false), (a => 253, b => 254, p => false), (a => 275, b => 276, p => false), (a => 297, b => 298, p => false), (a => 319, b => 320, p => false), (a => 341, b => 342, p => false), (a => 13, b => 14, p => false), (a => 35, b => 36, p => false), (a => 57, b => 58, p => false), (a => 79, b => 80, p => false), (a => 101, b => 102, p => false), (a => 123, b => 124, p => false), (a => 145, b => 146, p => false), (a => 167, b => 168, p => false), (a => 189, b => 190, p => false), (a => 211, b => 212, p => false), (a => 233, b => 234, p => false), (a => 255, b => 256, p => false), (a => 277, b => 278, p => false), (a => 299, b => 300, p => false), (a => 321, b => 322, p => false), (a => 343, b => 344, p => false), (a => 15, b => 16, p => false), (a => 37, b => 38, p => false), (a => 59, b => 60, p => false), (a => 81, b => 82, p => false), (a => 103, b => 104, p => false), (a => 125, b => 126, p => false), (a => 147, b => 148, p => false), (a => 169, b => 170, p => false), (a => 191, b => 192, p => false), (a => 213, b => 214, p => false), (a => 235, b => 236, p => false), (a => 257, b => 258, p => false), (a => 279, b => 280, p => false), (a => 301, b => 302, p => false), (a => 323, b => 324, p => false), (a => 345, b => 346, p => false), (a => 2, b => 24, p => false), (a => 46, b => 68, p => false), (a => 90, b => 112, p => false), (a => 134, b => 156, p => false), (a => 178, b => 200, p => false), (a => 222, b => 244, p => false), (a => 266, b => 288, p => false), (a => 310, b => 332, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 331, p => true), (a => 21, b => 330, p => true), (a => 22, b => 329, p => true), (a => 23, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 309, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 45, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 287, p => true), (a => 65, b => 286, p => true), (a => 66, b => 285, p => true), (a => 67, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 243, p => true), (a => 109, b => 242, p => true), (a => 110, b => 241, p => true), (a => 111, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 221, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 133, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 199, p => true), (a => 153, b => 198, p => true), (a => 154, b => 197, p => true), (a => 155, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 4, b => 5, p => false), (a => 26, b => 27, p => false), (a => 48, b => 49, p => false), (a => 70, b => 71, p => false), (a => 92, b => 93, p => false), (a => 114, b => 115, p => false), (a => 136, b => 137, p => false), (a => 158, b => 159, p => false), (a => 180, b => 181, p => false), (a => 202, b => 203, p => false), (a => 224, b => 225, p => false), (a => 246, b => 247, p => false), (a => 268, b => 269, p => false), (a => 290, b => 291, p => false), (a => 312, b => 313, p => false), (a => 334, b => 335, p => false), (a => 6, b => 7, p => false), (a => 28, b => 29, p => false), (a => 50, b => 51, p => false), (a => 72, b => 73, p => false), (a => 94, b => 95, p => false), (a => 116, b => 117, p => false), (a => 138, b => 139, p => false), (a => 160, b => 161, p => false), (a => 182, b => 183, p => false), (a => 204, b => 205, p => false), (a => 226, b => 227, p => false), (a => 248, b => 249, p => false), (a => 270, b => 271, p => false), (a => 292, b => 293, p => false), (a => 314, b => 315, p => false), (a => 336, b => 337, p => false), (a => 8, b => 9, p => false), (a => 30, b => 31, p => false), (a => 52, b => 53, p => false), (a => 74, b => 75, p => false), (a => 96, b => 97, p => false), (a => 118, b => 119, p => false), (a => 140, b => 141, p => false), (a => 162, b => 163, p => false), (a => 184, b => 185, p => false), (a => 206, b => 207, p => false), (a => 228, b => 229, p => false), (a => 250, b => 251, p => false), (a => 272, b => 273, p => false), (a => 294, b => 295, p => false), (a => 316, b => 317, p => false), (a => 338, b => 339, p => false), (a => 10, b => 11, p => false), (a => 32, b => 33, p => false), (a => 54, b => 55, p => false), (a => 76, b => 77, p => false), (a => 98, b => 99, p => false), (a => 120, b => 121, p => false), (a => 142, b => 143, p => false), (a => 164, b => 165, p => false), (a => 186, b => 187, p => false), (a => 208, b => 209, p => false), (a => 230, b => 231, p => false), (a => 252, b => 253, p => false), (a => 274, b => 275, p => false), (a => 296, b => 297, p => false), (a => 318, b => 319, p => false), (a => 340, b => 341, p => false), (a => 12, b => 13, p => false), (a => 34, b => 35, p => false), (a => 56, b => 57, p => false), (a => 78, b => 79, p => false), (a => 100, b => 101, p => false), (a => 122, b => 123, p => false), (a => 144, b => 145, p => false), (a => 166, b => 167, p => false), (a => 188, b => 189, p => false), (a => 210, b => 211, p => false), (a => 232, b => 233, p => false), (a => 254, b => 255, p => false), (a => 276, b => 277, p => false), (a => 298, b => 299, p => false), (a => 320, b => 321, p => false), (a => 342, b => 343, p => false), (a => 14, b => 15, p => false), (a => 36, b => 37, p => false), (a => 58, b => 59, p => false), (a => 80, b => 81, p => false), (a => 102, b => 103, p => false), (a => 124, b => 125, p => false), (a => 146, b => 147, p => false), (a => 168, b => 169, p => false), (a => 190, b => 191, p => false), (a => 212, b => 213, p => false), (a => 234, b => 235, p => false), (a => 256, b => 257, p => false), (a => 278, b => 279, p => false), (a => 300, b => 301, p => false), (a => 322, b => 323, p => false), (a => 344, b => 345, p => false), (a => 3, b => 25, p => false), (a => 47, b => 69, p => false), (a => 91, b => 113, p => false), (a => 135, b => 157, p => false), (a => 179, b => 201, p => false), (a => 223, b => 245, p => false), (a => 267, b => 289, p => false), (a => 311, b => 333, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 16, b => 348, p => true), (a => 17, b => 347, p => true), (a => 18, b => 346, p => true), (a => 19, b => 332, p => true), (a => 20, b => 331, p => true), (a => 21, b => 330, p => true), (a => 22, b => 329, p => true), (a => 23, b => 328, p => true), (a => 24, b => 327, p => true), (a => 38, b => 326, p => true), (a => 39, b => 325, p => true), (a => 40, b => 324, p => true), (a => 41, b => 310, p => true), (a => 42, b => 309, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 45, b => 306, p => true), (a => 46, b => 305, p => true), (a => 60, b => 304, p => true), (a => 61, b => 303, p => true), (a => 62, b => 302, p => true), (a => 63, b => 288, p => true), (a => 64, b => 287, p => true), (a => 65, b => 286, p => true), (a => 66, b => 285, p => true), (a => 67, b => 284, p => true), (a => 68, b => 283, p => true), (a => 82, b => 282, p => true), (a => 83, b => 281, p => true), (a => 84, b => 280, p => true), (a => 85, b => 266, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 90, b => 261, p => true), (a => 104, b => 260, p => true), (a => 105, b => 259, p => true), (a => 106, b => 258, p => true), (a => 107, b => 244, p => true), (a => 108, b => 243, p => true), (a => 109, b => 242, p => true), (a => 110, b => 241, p => true), (a => 111, b => 240, p => true), (a => 112, b => 239, p => true), (a => 126, b => 238, p => true), (a => 127, b => 237, p => true), (a => 128, b => 236, p => true), (a => 129, b => 222, p => true), (a => 130, b => 221, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 133, b => 218, p => true), (a => 134, b => 217, p => true), (a => 148, b => 216, p => true), (a => 149, b => 215, p => true), (a => 150, b => 214, p => true), (a => 151, b => 200, p => true), (a => 152, b => 199, p => true), (a => 153, b => 198, p => true), (a => 154, b => 197, p => true), (a => 155, b => 196, p => true), (a => 156, b => 195, p => true), (a => 170, b => 194, p => true), (a => 171, b => 193, p => true), (a => 172, b => 192, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 30, p => false), (a => 52, b => 74, p => false), (a => 96, b => 118, p => false), (a => 140, b => 162, p => false), (a => 184, b => 206, p => false), (a => 228, b => 250, p => false), (a => 272, b => 294, p => false), (a => 316, b => 338, p => false), (a => 4, b => 26, p => false), (a => 48, b => 70, p => false), (a => 92, b => 114, p => false), (a => 136, b => 158, p => false), (a => 180, b => 202, p => false), (a => 224, b => 246, p => false), (a => 268, b => 290, p => false), (a => 312, b => 334, p => false), (a => 12, b => 34, p => false), (a => 56, b => 78, p => false), (a => 100, b => 122, p => false), (a => 144, b => 166, p => false), (a => 188, b => 210, p => false), (a => 232, b => 254, p => false), (a => 276, b => 298, p => false), (a => 320, b => 342, p => false), (a => 10, b => 32, p => false), (a => 54, b => 76, p => false), (a => 98, b => 120, p => false), (a => 142, b => 164, p => false), (a => 186, b => 208, p => false), (a => 230, b => 252, p => false), (a => 274, b => 296, p => false), (a => 318, b => 340, p => false), (a => 6, b => 28, p => false), (a => 50, b => 72, p => false), (a => 94, b => 116, p => false), (a => 138, b => 160, p => false), (a => 182, b => 204, p => false), (a => 226, b => 248, p => false), (a => 270, b => 292, p => false), (a => 314, b => 336, p => false), (a => 14, b => 36, p => false), (a => 58, b => 80, p => false), (a => 102, b => 124, p => false), (a => 146, b => 168, p => false), (a => 190, b => 212, p => false), (a => 234, b => 256, p => false), (a => 278, b => 300, p => false), (a => 322, b => 344, p => false), (a => 9, b => 31, p => false), (a => 53, b => 75, p => false), (a => 97, b => 119, p => false), (a => 141, b => 163, p => false), (a => 185, b => 207, p => false), (a => 229, b => 251, p => false), (a => 273, b => 295, p => false), (a => 317, b => 339, p => false), (a => 5, b => 27, p => false), (a => 49, b => 71, p => false), (a => 93, b => 115, p => false), (a => 137, b => 159, p => false), (a => 181, b => 203, p => false), (a => 225, b => 247, p => false), (a => 269, b => 291, p => false), (a => 313, b => 335, p => false), (a => 13, b => 35, p => false), (a => 57, b => 79, p => false), (a => 101, b => 123, p => false), (a => 145, b => 167, p => false), (a => 189, b => 211, p => false), (a => 233, b => 255, p => false), (a => 277, b => 299, p => false), (a => 321, b => 343, p => false), (a => 11, b => 33, p => false), (a => 55, b => 77, p => false), (a => 99, b => 121, p => false), (a => 143, b => 165, p => false), (a => 187, b => 209, p => false), (a => 231, b => 253, p => false), (a => 275, b => 297, p => false), (a => 319, b => 341, p => false), (a => 7, b => 29, p => false), (a => 51, b => 73, p => false), (a => 95, b => 117, p => false), (a => 139, b => 161, p => false), (a => 183, b => 205, p => false), (a => 227, b => 249, p => false), (a => 271, b => 293, p => false), (a => 315, b => 337, p => false), (a => 15, b => 37, p => false), (a => 59, b => 81, p => false), (a => 103, b => 125, p => false), (a => 147, b => 169, p => false), (a => 191, b => 213, p => false), (a => 235, b => 257, p => false), (a => 279, b => 301, p => false), (a => 323, b => 345, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 16, b => 347, p => true), (a => 17, b => 346, p => true), (a => 18, b => 333, p => true), (a => 19, b => 332, p => true), (a => 20, b => 331, p => true), (a => 21, b => 330, p => true), (a => 22, b => 329, p => true), (a => 23, b => 328, p => true), (a => 24, b => 327, p => true), (a => 25, b => 326, p => true), (a => 38, b => 325, p => true), (a => 39, b => 324, p => true), (a => 40, b => 311, p => true), (a => 41, b => 310, p => true), (a => 42, b => 309, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 45, b => 306, p => true), (a => 46, b => 305, p => true), (a => 47, b => 304, p => true), (a => 60, b => 303, p => true), (a => 61, b => 302, p => true), (a => 62, b => 289, p => true), (a => 63, b => 288, p => true), (a => 64, b => 287, p => true), (a => 65, b => 286, p => true), (a => 66, b => 285, p => true), (a => 67, b => 284, p => true), (a => 68, b => 283, p => true), (a => 69, b => 282, p => true), (a => 82, b => 281, p => true), (a => 83, b => 280, p => true), (a => 84, b => 267, p => true), (a => 85, b => 266, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 90, b => 261, p => true), (a => 91, b => 260, p => true), (a => 104, b => 259, p => true), (a => 105, b => 258, p => true), (a => 106, b => 245, p => true), (a => 107, b => 244, p => true), (a => 108, b => 243, p => true), (a => 109, b => 242, p => true), (a => 110, b => 241, p => true), (a => 111, b => 240, p => true), (a => 112, b => 239, p => true), (a => 113, b => 238, p => true), (a => 126, b => 237, p => true), (a => 127, b => 236, p => true), (a => 128, b => 223, p => true), (a => 129, b => 222, p => true), (a => 130, b => 221, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 133, b => 218, p => true), (a => 134, b => 217, p => true), (a => 135, b => 216, p => true), (a => 148, b => 215, p => true), (a => 149, b => 214, p => true), (a => 150, b => 201, p => true), (a => 151, b => 200, p => true), (a => 152, b => 199, p => true), (a => 153, b => 198, p => true), (a => 154, b => 197, p => true), (a => 155, b => 196, p => true), (a => 156, b => 195, p => true), (a => 157, b => 194, p => true), (a => 170, b => 193, p => true), (a => 171, b => 192, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 22, p => false), (a => 52, b => 66, p => false), (a => 96, b => 110, p => false), (a => 140, b => 154, p => false), (a => 184, b => 198, p => false), (a => 228, b => 242, p => false), (a => 272, b => 286, p => false), (a => 316, b => 330, p => false), (a => 12, b => 26, p => false), (a => 56, b => 70, p => false), (a => 100, b => 114, p => false), (a => 144, b => 158, p => false), (a => 188, b => 202, p => false), (a => 232, b => 246, p => false), (a => 276, b => 290, p => false), (a => 320, b => 334, p => false), (a => 10, b => 24, p => false), (a => 54, b => 68, p => false), (a => 98, b => 112, p => false), (a => 142, b => 156, p => false), (a => 186, b => 200, p => false), (a => 230, b => 244, p => false), (a => 274, b => 288, p => false), (a => 318, b => 332, p => false), (a => 14, b => 28, p => false), (a => 58, b => 72, p => false), (a => 102, b => 116, p => false), (a => 146, b => 160, p => false), (a => 190, b => 204, p => false), (a => 234, b => 248, p => false), (a => 278, b => 292, p => false), (a => 322, b => 336, p => false), (a => 9, b => 23, p => false), (a => 53, b => 67, p => false), (a => 97, b => 111, p => false), (a => 141, b => 155, p => false), (a => 185, b => 199, p => false), (a => 229, b => 243, p => false), (a => 273, b => 287, p => false), (a => 317, b => 331, p => false), (a => 13, b => 27, p => false), (a => 57, b => 71, p => false), (a => 101, b => 115, p => false), (a => 145, b => 159, p => false), (a => 189, b => 203, p => false), (a => 233, b => 247, p => false), (a => 277, b => 291, p => false), (a => 321, b => 335, p => false), (a => 11, b => 25, p => false), (a => 55, b => 69, p => false), (a => 99, b => 113, p => false), (a => 143, b => 157, p => false), (a => 187, b => 201, p => false), (a => 231, b => 245, p => false), (a => 275, b => 289, p => false), (a => 319, b => 333, p => false), (a => 15, b => 29, p => false), (a => 59, b => 73, p => false), (a => 103, b => 117, p => false), (a => 147, b => 161, p => false), (a => 191, b => 205, p => false), (a => 235, b => 249, p => false), (a => 279, b => 293, p => false), (a => 323, b => 337, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 4, b => 347, p => true), (a => 5, b => 346, p => true), (a => 6, b => 345, p => true), (a => 7, b => 344, p => true), (a => 16, b => 343, p => true), (a => 17, b => 342, p => true), (a => 18, b => 341, p => true), (a => 19, b => 340, p => true), (a => 20, b => 339, p => true), (a => 21, b => 338, p => true), (a => 30, b => 329, p => true), (a => 31, b => 328, p => true), (a => 32, b => 327, p => true), (a => 33, b => 326, p => true), (a => 34, b => 325, p => true), (a => 35, b => 324, p => true), (a => 36, b => 315, p => true), (a => 37, b => 314, p => true), (a => 38, b => 313, p => true), (a => 39, b => 312, p => true), (a => 40, b => 311, p => true), (a => 41, b => 310, p => true), (a => 42, b => 309, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 45, b => 306, p => true), (a => 46, b => 305, p => true), (a => 47, b => 304, p => true), (a => 48, b => 303, p => true), (a => 49, b => 302, p => true), (a => 50, b => 301, p => true), (a => 51, b => 300, p => true), (a => 60, b => 299, p => true), (a => 61, b => 298, p => true), (a => 62, b => 297, p => true), (a => 63, b => 296, p => true), (a => 64, b => 295, p => true), (a => 65, b => 294, p => true), (a => 74, b => 285, p => true), (a => 75, b => 284, p => true), (a => 76, b => 283, p => true), (a => 77, b => 282, p => true), (a => 78, b => 281, p => true), (a => 79, b => 280, p => true), (a => 80, b => 271, p => true), (a => 81, b => 270, p => true), (a => 82, b => 269, p => true), (a => 83, b => 268, p => true), (a => 84, b => 267, p => true), (a => 85, b => 266, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 90, b => 261, p => true), (a => 91, b => 260, p => true), (a => 92, b => 259, p => true), (a => 93, b => 258, p => true), (a => 94, b => 257, p => true), (a => 95, b => 256, p => true), (a => 104, b => 255, p => true), (a => 105, b => 254, p => true), (a => 106, b => 253, p => true), (a => 107, b => 252, p => true), (a => 108, b => 251, p => true), (a => 109, b => 250, p => true), (a => 118, b => 241, p => true), (a => 119, b => 240, p => true), (a => 120, b => 239, p => true), (a => 121, b => 238, p => true), (a => 122, b => 237, p => true), (a => 123, b => 236, p => true), (a => 124, b => 227, p => true), (a => 125, b => 226, p => true), (a => 126, b => 225, p => true), (a => 127, b => 224, p => true), (a => 128, b => 223, p => true), (a => 129, b => 222, p => true), (a => 130, b => 221, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 133, b => 218, p => true), (a => 134, b => 217, p => true), (a => 135, b => 216, p => true), (a => 136, b => 215, p => true), (a => 137, b => 214, p => true), (a => 138, b => 213, p => true), (a => 139, b => 212, p => true), (a => 148, b => 211, p => true), (a => 149, b => 210, p => true), (a => 150, b => 209, p => true), (a => 151, b => 208, p => true), (a => 152, b => 207, p => true), (a => 153, b => 206, p => true), (a => 162, b => 197, p => true), (a => 163, b => 196, p => true), (a => 164, b => 195, p => true), (a => 165, b => 194, p => true), (a => 166, b => 193, p => true), (a => 167, b => 192, p => true), (a => 168, b => 183, p => true), (a => 169, b => 182, p => true), (a => 170, b => 181, p => true), (a => 171, b => 180, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 4, b => 8, p => false), (a => 48, b => 52, p => false), (a => 92, b => 96, p => false), (a => 136, b => 140, p => false), (a => 180, b => 184, p => false), (a => 224, b => 228, p => false), (a => 268, b => 272, p => false), (a => 312, b => 316, p => false), (a => 12, b => 22, p => false), (a => 56, b => 66, p => false), (a => 100, b => 110, p => false), (a => 144, b => 154, p => false), (a => 188, b => 198, p => false), (a => 232, b => 242, p => false), (a => 276, b => 286, p => false), (a => 320, b => 330, p => false), (a => 6, b => 10, p => false), (a => 50, b => 54, p => false), (a => 94, b => 98, p => false), (a => 138, b => 142, p => false), (a => 182, b => 186, p => false), (a => 226, b => 230, p => false), (a => 270, b => 274, p => false), (a => 314, b => 318, p => false), (a => 14, b => 24, p => false), (a => 58, b => 68, p => false), (a => 102, b => 112, p => false), (a => 146, b => 156, p => false), (a => 190, b => 200, p => false), (a => 234, b => 244, p => false), (a => 278, b => 288, p => false), (a => 322, b => 332, p => false), (a => 5, b => 9, p => false), (a => 49, b => 53, p => false), (a => 93, b => 97, p => false), (a => 137, b => 141, p => false), (a => 181, b => 185, p => false), (a => 225, b => 229, p => false), (a => 269, b => 273, p => false), (a => 313, b => 317, p => false), (a => 13, b => 23, p => false), (a => 57, b => 67, p => false), (a => 101, b => 111, p => false), (a => 145, b => 155, p => false), (a => 189, b => 199, p => false), (a => 233, b => 243, p => false), (a => 277, b => 287, p => false), (a => 321, b => 331, p => false), (a => 7, b => 11, p => false), (a => 51, b => 55, p => false), (a => 95, b => 99, p => false), (a => 139, b => 143, p => false), (a => 183, b => 187, p => false), (a => 227, b => 231, p => false), (a => 271, b => 275, p => false), (a => 315, b => 319, p => false), (a => 15, b => 25, p => false), (a => 59, b => 69, p => false), (a => 103, b => 113, p => false), (a => 147, b => 157, p => false), (a => 191, b => 201, p => false), (a => 235, b => 245, p => false), (a => 279, b => 289, p => false), (a => 323, b => 333, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 16, b => 347, p => true), (a => 17, b => 346, p => true), (a => 18, b => 345, p => true), (a => 19, b => 344, p => true), (a => 20, b => 343, p => true), (a => 21, b => 342, p => true), (a => 26, b => 341, p => true), (a => 27, b => 340, p => true), (a => 28, b => 339, p => true), (a => 29, b => 338, p => true), (a => 30, b => 337, p => true), (a => 31, b => 336, p => true), (a => 32, b => 335, p => true), (a => 33, b => 334, p => true), (a => 34, b => 329, p => true), (a => 35, b => 328, p => true), (a => 36, b => 327, p => true), (a => 37, b => 326, p => true), (a => 38, b => 325, p => true), (a => 39, b => 324, p => true), (a => 40, b => 311, p => true), (a => 41, b => 310, p => true), (a => 42, b => 309, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 45, b => 306, p => true), (a => 46, b => 305, p => true), (a => 47, b => 304, p => true), (a => 60, b => 303, p => true), (a => 61, b => 302, p => true), (a => 62, b => 301, p => true), (a => 63, b => 300, p => true), (a => 64, b => 299, p => true), (a => 65, b => 298, p => true), (a => 70, b => 297, p => true), (a => 71, b => 296, p => true), (a => 72, b => 295, p => true), (a => 73, b => 294, p => true), (a => 74, b => 293, p => true), (a => 75, b => 292, p => true), (a => 76, b => 291, p => true), (a => 77, b => 290, p => true), (a => 78, b => 285, p => true), (a => 79, b => 284, p => true), (a => 80, b => 283, p => true), (a => 81, b => 282, p => true), (a => 82, b => 281, p => true), (a => 83, b => 280, p => true), (a => 84, b => 267, p => true), (a => 85, b => 266, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 90, b => 261, p => true), (a => 91, b => 260, p => true), (a => 104, b => 259, p => true), (a => 105, b => 258, p => true), (a => 106, b => 257, p => true), (a => 107, b => 256, p => true), (a => 108, b => 255, p => true), (a => 109, b => 254, p => true), (a => 114, b => 253, p => true), (a => 115, b => 252, p => true), (a => 116, b => 251, p => true), (a => 117, b => 250, p => true), (a => 118, b => 249, p => true), (a => 119, b => 248, p => true), (a => 120, b => 247, p => true), (a => 121, b => 246, p => true), (a => 122, b => 241, p => true), (a => 123, b => 240, p => true), (a => 124, b => 239, p => true), (a => 125, b => 238, p => true), (a => 126, b => 237, p => true), (a => 127, b => 236, p => true), (a => 128, b => 223, p => true), (a => 129, b => 222, p => true), (a => 130, b => 221, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 133, b => 218, p => true), (a => 134, b => 217, p => true), (a => 135, b => 216, p => true), (a => 148, b => 215, p => true), (a => 149, b => 214, p => true), (a => 150, b => 213, p => true), (a => 151, b => 212, p => true), (a => 152, b => 211, p => true), (a => 153, b => 210, p => true), (a => 158, b => 209, p => true), (a => 159, b => 208, p => true), (a => 160, b => 207, p => true), (a => 161, b => 206, p => true), (a => 162, b => 205, p => true), (a => 163, b => 204, p => true), (a => 164, b => 203, p => true), (a => 165, b => 202, p => true), (a => 166, b => 197, p => true), (a => 167, b => 196, p => true), (a => 168, b => 195, p => true), (a => 169, b => 194, p => true), (a => 170, b => 193, p => true), (a => 171, b => 192, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 2, b => 4, p => false), (a => 46, b => 48, p => false), (a => 90, b => 92, p => false), (a => 134, b => 136, p => false), (a => 178, b => 180, p => false), (a => 222, b => 224, p => false), (a => 266, b => 268, p => false), (a => 310, b => 312, p => false), (a => 6, b => 8, p => false), (a => 50, b => 52, p => false), (a => 94, b => 96, p => false), (a => 138, b => 140, p => false), (a => 182, b => 184, p => false), (a => 226, b => 228, p => false), (a => 270, b => 272, p => false), (a => 314, b => 316, p => false), (a => 10, b => 12, p => false), (a => 54, b => 56, p => false), (a => 98, b => 100, p => false), (a => 142, b => 144, p => false), (a => 186, b => 188, p => false), (a => 230, b => 232, p => false), (a => 274, b => 276, p => false), (a => 318, b => 320, p => false), (a => 14, b => 22, p => false), (a => 58, b => 66, p => false), (a => 102, b => 110, p => false), (a => 146, b => 154, p => false), (a => 190, b => 198, p => false), (a => 234, b => 242, p => false), (a => 278, b => 286, p => false), (a => 322, b => 330, p => false), (a => 3, b => 5, p => false), (a => 47, b => 49, p => false), (a => 91, b => 93, p => false), (a => 135, b => 137, p => false), (a => 179, b => 181, p => false), (a => 223, b => 225, p => false), (a => 267, b => 269, p => false), (a => 311, b => 313, p => false), (a => 7, b => 9, p => false), (a => 51, b => 53, p => false), (a => 95, b => 97, p => false), (a => 139, b => 141, p => false), (a => 183, b => 185, p => false), (a => 227, b => 229, p => false), (a => 271, b => 273, p => false), (a => 315, b => 317, p => false), (a => 11, b => 13, p => false), (a => 55, b => 57, p => false), (a => 99, b => 101, p => false), (a => 143, b => 145, p => false), (a => 187, b => 189, p => false), (a => 231, b => 233, p => false), (a => 275, b => 277, p => false), (a => 319, b => 321, p => false), (a => 15, b => 23, p => false), (a => 59, b => 67, p => false), (a => 103, b => 111, p => false), (a => 147, b => 155, p => false), (a => 191, b => 199, p => false), (a => 235, b => 243, p => false), (a => 279, b => 287, p => false), (a => 323, b => 331, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 16, b => 349, p => true), (a => 17, b => 348, p => true), (a => 18, b => 347, p => true), (a => 19, b => 346, p => true), (a => 20, b => 345, p => true), (a => 21, b => 344, p => true), (a => 24, b => 343, p => true), (a => 25, b => 342, p => true), (a => 26, b => 341, p => true), (a => 27, b => 340, p => true), (a => 28, b => 339, p => true), (a => 29, b => 338, p => true), (a => 30, b => 337, p => true), (a => 31, b => 336, p => true), (a => 32, b => 335, p => true), (a => 33, b => 334, p => true), (a => 34, b => 333, p => true), (a => 35, b => 332, p => true), (a => 36, b => 329, p => true), (a => 37, b => 328, p => true), (a => 38, b => 327, p => true), (a => 39, b => 326, p => true), (a => 40, b => 325, p => true), (a => 41, b => 324, p => true), (a => 42, b => 309, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 45, b => 306, p => true), (a => 60, b => 305, p => true), (a => 61, b => 304, p => true), (a => 62, b => 303, p => true), (a => 63, b => 302, p => true), (a => 64, b => 301, p => true), (a => 65, b => 300, p => true), (a => 68, b => 299, p => true), (a => 69, b => 298, p => true), (a => 70, b => 297, p => true), (a => 71, b => 296, p => true), (a => 72, b => 295, p => true), (a => 73, b => 294, p => true), (a => 74, b => 293, p => true), (a => 75, b => 292, p => true), (a => 76, b => 291, p => true), (a => 77, b => 290, p => true), (a => 78, b => 289, p => true), (a => 79, b => 288, p => true), (a => 80, b => 285, p => true), (a => 81, b => 284, p => true), (a => 82, b => 283, p => true), (a => 83, b => 282, p => true), (a => 84, b => 281, p => true), (a => 85, b => 280, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 104, b => 261, p => true), (a => 105, b => 260, p => true), (a => 106, b => 259, p => true), (a => 107, b => 258, p => true), (a => 108, b => 257, p => true), (a => 109, b => 256, p => true), (a => 112, b => 255, p => true), (a => 113, b => 254, p => true), (a => 114, b => 253, p => true), (a => 115, b => 252, p => true), (a => 116, b => 251, p => true), (a => 117, b => 250, p => true), (a => 118, b => 249, p => true), (a => 119, b => 248, p => true), (a => 120, b => 247, p => true), (a => 121, b => 246, p => true), (a => 122, b => 245, p => true), (a => 123, b => 244, p => true), (a => 124, b => 241, p => true), (a => 125, b => 240, p => true), (a => 126, b => 239, p => true), (a => 127, b => 238, p => true), (a => 128, b => 237, p => true), (a => 129, b => 236, p => true), (a => 130, b => 221, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 133, b => 218, p => true), (a => 148, b => 217, p => true), (a => 149, b => 216, p => true), (a => 150, b => 215, p => true), (a => 151, b => 214, p => true), (a => 152, b => 213, p => true), (a => 153, b => 212, p => true), (a => 156, b => 211, p => true), (a => 157, b => 210, p => true), (a => 158, b => 209, p => true), (a => 159, b => 208, p => true), (a => 160, b => 207, p => true), (a => 161, b => 206, p => true), (a => 162, b => 205, p => true), (a => 163, b => 204, p => true), (a => 164, b => 203, p => true), (a => 165, b => 202, p => true), (a => 166, b => 201, p => true), (a => 167, b => 200, p => true), (a => 168, b => 197, p => true), (a => 169, b => 196, p => true), (a => 170, b => 195, p => true), (a => 171, b => 194, p => true), (a => 172, b => 193, p => true), (a => 173, b => 192, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 1, b => 2, p => false), (a => 45, b => 46, p => false), (a => 89, b => 90, p => false), (a => 133, b => 134, p => false), (a => 177, b => 178, p => false), (a => 221, b => 222, p => false), (a => 265, b => 266, p => false), (a => 309, b => 310, p => false), (a => 3, b => 4, p => false), (a => 47, b => 48, p => false), (a => 91, b => 92, p => false), (a => 135, b => 136, p => false), (a => 179, b => 180, p => false), (a => 223, b => 224, p => false), (a => 267, b => 268, p => false), (a => 311, b => 312, p => false), (a => 5, b => 6, p => false), (a => 49, b => 50, p => false), (a => 93, b => 94, p => false), (a => 137, b => 138, p => false), (a => 181, b => 182, p => false), (a => 225, b => 226, p => false), (a => 269, b => 270, p => false), (a => 313, b => 314, p => false), (a => 7, b => 8, p => false), (a => 51, b => 52, p => false), (a => 95, b => 96, p => false), (a => 139, b => 140, p => false), (a => 183, b => 184, p => false), (a => 227, b => 228, p => false), (a => 271, b => 272, p => false), (a => 315, b => 316, p => false), (a => 9, b => 10, p => false), (a => 53, b => 54, p => false), (a => 97, b => 98, p => false), (a => 141, b => 142, p => false), (a => 185, b => 186, p => false), (a => 229, b => 230, p => false), (a => 273, b => 274, p => false), (a => 317, b => 318, p => false), (a => 11, b => 12, p => false), (a => 55, b => 56, p => false), (a => 99, b => 100, p => false), (a => 143, b => 144, p => false), (a => 187, b => 188, p => false), (a => 231, b => 232, p => false), (a => 275, b => 276, p => false), (a => 319, b => 320, p => false), (a => 13, b => 14, p => false), (a => 57, b => 58, p => false), (a => 101, b => 102, p => false), (a => 145, b => 146, p => false), (a => 189, b => 190, p => false), (a => 233, b => 234, p => false), (a => 277, b => 278, p => false), (a => 321, b => 322, p => false), (a => 15, b => 22, p => false), (a => 59, b => 66, p => false), (a => 103, b => 110, p => false), (a => 147, b => 154, p => false), (a => 191, b => 198, p => false), (a => 235, b => 242, p => false), (a => 279, b => 286, p => false), (a => 323, b => 330, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 23, b => 344, p => true), (a => 24, b => 343, p => true), (a => 25, b => 342, p => true), (a => 26, b => 341, p => true), (a => 27, b => 340, p => true), (a => 28, b => 339, p => true), (a => 29, b => 338, p => true), (a => 30, b => 337, p => true), (a => 31, b => 336, p => true), (a => 32, b => 335, p => true), (a => 33, b => 334, p => true), (a => 34, b => 333, p => true), (a => 35, b => 332, p => true), (a => 36, b => 331, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 67, b => 300, p => true), (a => 68, b => 299, p => true), (a => 69, b => 298, p => true), (a => 70, b => 297, p => true), (a => 71, b => 296, p => true), (a => 72, b => 295, p => true), (a => 73, b => 294, p => true), (a => 74, b => 293, p => true), (a => 75, b => 292, p => true), (a => 76, b => 291, p => true), (a => 77, b => 290, p => true), (a => 78, b => 289, p => true), (a => 79, b => 288, p => true), (a => 80, b => 287, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 111, b => 256, p => true), (a => 112, b => 255, p => true), (a => 113, b => 254, p => true), (a => 114, b => 253, p => true), (a => 115, b => 252, p => true), (a => 116, b => 251, p => true), (a => 117, b => 250, p => true), (a => 118, b => 249, p => true), (a => 119, b => 248, p => true), (a => 120, b => 247, p => true), (a => 121, b => 246, p => true), (a => 122, b => 245, p => true), (a => 123, b => 244, p => true), (a => 124, b => 243, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 155, b => 212, p => true), (a => 156, b => 211, p => true), (a => 157, b => 210, p => true), (a => 158, b => 209, p => true), (a => 159, b => 208, p => true), (a => 160, b => 207, p => true), (a => 161, b => 206, p => true), (a => 162, b => 205, p => true), (a => 163, b => 204, p => true), (a => 164, b => 203, p => true), (a => 165, b => 202, p => true), (a => 166, b => 201, p => true), (a => 167, b => 200, p => true), (a => 168, b => 199, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 52, p => false), (a => 96, b => 140, p => false), (a => 184, b => 228, p => false), (a => 272, b => 316, p => false), (a => 4, b => 48, p => false), (a => 92, b => 136, p => false), (a => 180, b => 224, p => false), (a => 268, b => 312, p => false), (a => 12, b => 56, p => false), (a => 100, b => 144, p => false), (a => 188, b => 232, p => false), (a => 276, b => 320, p => false), (a => 2, b => 46, p => false), (a => 90, b => 134, p => false), (a => 178, b => 222, p => false), (a => 266, b => 310, p => false), (a => 10, b => 54, p => false), (a => 98, b => 142, p => false), (a => 186, b => 230, p => false), (a => 274, b => 318, p => false), (a => 6, b => 50, p => false), (a => 94, b => 138, p => false), (a => 182, b => 226, p => false), (a => 270, b => 314, p => false), (a => 14, b => 58, p => false), (a => 102, b => 146, p => false), (a => 190, b => 234, p => false), (a => 278, b => 322, p => false), (a => 1, b => 45, p => false), (a => 89, b => 133, p => false), (a => 177, b => 221, p => false), (a => 265, b => 309, p => false), (a => 9, b => 53, p => false), (a => 97, b => 141, p => false), (a => 185, b => 229, p => false), (a => 273, b => 317, p => false), (a => 5, b => 49, p => false), (a => 93, b => 137, p => false), (a => 181, b => 225, p => false), (a => 269, b => 313, p => false), (a => 13, b => 57, p => false), (a => 101, b => 145, p => false), (a => 189, b => 233, p => false), (a => 277, b => 321, p => false), (a => 3, b => 47, p => false), (a => 91, b => 135, p => false), (a => 179, b => 223, p => false), (a => 267, b => 311, p => false), (a => 11, b => 55, p => false), (a => 99, b => 143, p => false), (a => 187, b => 231, p => false), (a => 275, b => 319, p => false), (a => 7, b => 51, p => false), (a => 95, b => 139, p => false), (a => 183, b => 227, p => false), (a => 271, b => 315, p => false), (a => 15, b => 59, p => false), (a => 103, b => 147, p => false), (a => 191, b => 235, p => false), (a => 279, b => 323, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 22, b => 344, p => true), (a => 23, b => 343, p => true), (a => 24, b => 342, p => true), (a => 25, b => 341, p => true), (a => 26, b => 340, p => true), (a => 27, b => 339, p => true), (a => 28, b => 338, p => true), (a => 29, b => 337, p => true), (a => 30, b => 336, p => true), (a => 31, b => 335, p => true), (a => 32, b => 334, p => true), (a => 33, b => 333, p => true), (a => 34, b => 332, p => true), (a => 35, b => 331, p => true), (a => 36, b => 330, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 308, p => true), (a => 44, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 66, b => 300, p => true), (a => 67, b => 299, p => true), (a => 68, b => 298, p => true), (a => 69, b => 297, p => true), (a => 70, b => 296, p => true), (a => 71, b => 295, p => true), (a => 72, b => 294, p => true), (a => 73, b => 293, p => true), (a => 74, b => 292, p => true), (a => 75, b => 291, p => true), (a => 76, b => 290, p => true), (a => 77, b => 289, p => true), (a => 78, b => 288, p => true), (a => 79, b => 287, p => true), (a => 80, b => 286, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 110, b => 256, p => true), (a => 111, b => 255, p => true), (a => 112, b => 254, p => true), (a => 113, b => 253, p => true), (a => 114, b => 252, p => true), (a => 115, b => 251, p => true), (a => 116, b => 250, p => true), (a => 117, b => 249, p => true), (a => 118, b => 248, p => true), (a => 119, b => 247, p => true), (a => 120, b => 246, p => true), (a => 121, b => 245, p => true), (a => 122, b => 244, p => true), (a => 123, b => 243, p => true), (a => 124, b => 242, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 220, p => true), (a => 132, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 154, b => 212, p => true), (a => 155, b => 211, p => true), (a => 156, b => 210, p => true), (a => 157, b => 209, p => true), (a => 158, b => 208, p => true), (a => 159, b => 207, p => true), (a => 160, b => 206, p => true), (a => 161, b => 205, p => true), (a => 162, b => 204, p => true), (a => 163, b => 203, p => true), (a => 164, b => 202, p => true), (a => 165, b => 201, p => true), (a => 166, b => 200, p => true), (a => 167, b => 199, p => true), (a => 168, b => 198, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 44, p => false), (a => 96, b => 132, p => false), (a => 184, b => 220, p => false), (a => 272, b => 308, p => false), (a => 12, b => 48, p => false), (a => 100, b => 136, p => false), (a => 188, b => 224, p => false), (a => 276, b => 312, p => false), (a => 10, b => 46, p => false), (a => 98, b => 134, p => false), (a => 186, b => 222, p => false), (a => 274, b => 310, p => false), (a => 14, b => 50, p => false), (a => 102, b => 138, p => false), (a => 190, b => 226, p => false), (a => 278, b => 314, p => false), (a => 9, b => 45, p => false), (a => 97, b => 133, p => false), (a => 185, b => 221, p => false), (a => 273, b => 309, p => false), (a => 13, b => 49, p => false), (a => 101, b => 137, p => false), (a => 189, b => 225, p => false), (a => 277, b => 313, p => false), (a => 11, b => 47, p => false), (a => 99, b => 135, p => false), (a => 187, b => 223, p => false), (a => 275, b => 311, p => false), (a => 15, b => 51, p => false), (a => 103, b => 139, p => false), (a => 191, b => 227, p => false), (a => 279, b => 315, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 4, b => 347, p => true), (a => 5, b => 346, p => true), (a => 6, b => 345, p => true), (a => 7, b => 344, p => true), (a => 16, b => 343, p => true), (a => 17, b => 342, p => true), (a => 18, b => 341, p => true), (a => 19, b => 340, p => true), (a => 20, b => 339, p => true), (a => 21, b => 338, p => true), (a => 22, b => 337, p => true), (a => 23, b => 336, p => true), (a => 24, b => 335, p => true), (a => 25, b => 334, p => true), (a => 26, b => 333, p => true), (a => 27, b => 332, p => true), (a => 28, b => 331, p => true), (a => 29, b => 330, p => true), (a => 30, b => 329, p => true), (a => 31, b => 328, p => true), (a => 32, b => 327, p => true), (a => 33, b => 326, p => true), (a => 34, b => 325, p => true), (a => 35, b => 324, p => true), (a => 36, b => 323, p => true), (a => 37, b => 322, p => true), (a => 38, b => 321, p => true), (a => 39, b => 320, p => true), (a => 40, b => 319, p => true), (a => 41, b => 318, p => true), (a => 42, b => 317, p => true), (a => 43, b => 316, p => true), (a => 52, b => 307, p => true), (a => 53, b => 306, p => true), (a => 54, b => 305, p => true), (a => 55, b => 304, p => true), (a => 56, b => 303, p => true), (a => 57, b => 302, p => true), (a => 58, b => 301, p => true), (a => 59, b => 300, p => true), (a => 60, b => 299, p => true), (a => 61, b => 298, p => true), (a => 62, b => 297, p => true), (a => 63, b => 296, p => true), (a => 64, b => 295, p => true), (a => 65, b => 294, p => true), (a => 66, b => 293, p => true), (a => 67, b => 292, p => true), (a => 68, b => 291, p => true), (a => 69, b => 290, p => true), (a => 70, b => 289, p => true), (a => 71, b => 288, p => true), (a => 72, b => 287, p => true), (a => 73, b => 286, p => true), (a => 74, b => 285, p => true), (a => 75, b => 284, p => true), (a => 76, b => 283, p => true), (a => 77, b => 282, p => true), (a => 78, b => 281, p => true), (a => 79, b => 280, p => true), (a => 80, b => 271, p => true), (a => 81, b => 270, p => true), (a => 82, b => 269, p => true), (a => 83, b => 268, p => true), (a => 84, b => 267, p => true), (a => 85, b => 266, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 90, b => 261, p => true), (a => 91, b => 260, p => true), (a => 92, b => 259, p => true), (a => 93, b => 258, p => true), (a => 94, b => 257, p => true), (a => 95, b => 256, p => true), (a => 104, b => 255, p => true), (a => 105, b => 254, p => true), (a => 106, b => 253, p => true), (a => 107, b => 252, p => true), (a => 108, b => 251, p => true), (a => 109, b => 250, p => true), (a => 110, b => 249, p => true), (a => 111, b => 248, p => true), (a => 112, b => 247, p => true), (a => 113, b => 246, p => true), (a => 114, b => 245, p => true), (a => 115, b => 244, p => true), (a => 116, b => 243, p => true), (a => 117, b => 242, p => true), (a => 118, b => 241, p => true), (a => 119, b => 240, p => true), (a => 120, b => 239, p => true), (a => 121, b => 238, p => true), (a => 122, b => 237, p => true), (a => 123, b => 236, p => true), (a => 124, b => 235, p => true), (a => 125, b => 234, p => true), (a => 126, b => 233, p => true), (a => 127, b => 232, p => true), (a => 128, b => 231, p => true), (a => 129, b => 230, p => true), (a => 130, b => 229, p => true), (a => 131, b => 228, p => true), (a => 140, b => 219, p => true), (a => 141, b => 218, p => true), (a => 142, b => 217, p => true), (a => 143, b => 216, p => true), (a => 144, b => 215, p => true), (a => 145, b => 214, p => true), (a => 146, b => 213, p => true), (a => 147, b => 212, p => true), (a => 148, b => 211, p => true), (a => 149, b => 210, p => true), (a => 150, b => 209, p => true), (a => 151, b => 208, p => true), (a => 152, b => 207, p => true), (a => 153, b => 206, p => true), (a => 154, b => 205, p => true), (a => 155, b => 204, p => true), (a => 156, b => 203, p => true), (a => 157, b => 202, p => true), (a => 158, b => 201, p => true), (a => 159, b => 200, p => true), (a => 160, b => 199, p => true), (a => 161, b => 198, p => true), (a => 162, b => 197, p => true), (a => 163, b => 196, p => true), (a => 164, b => 195, p => true), (a => 165, b => 194, p => true), (a => 166, b => 193, p => true), (a => 167, b => 192, p => true), (a => 168, b => 183, p => true), (a => 169, b => 182, p => true), (a => 170, b => 181, p => true), (a => 171, b => 180, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 4, b => 8, p => false), (a => 92, b => 96, p => false), (a => 180, b => 184, p => false), (a => 268, b => 272, p => false), (a => 12, b => 44, p => false), (a => 100, b => 132, p => false), (a => 188, b => 220, p => false), (a => 276, b => 308, p => false), (a => 6, b => 10, p => false), (a => 94, b => 98, p => false), (a => 182, b => 186, p => false), (a => 270, b => 274, p => false), (a => 14, b => 46, p => false), (a => 102, b => 134, p => false), (a => 190, b => 222, p => false), (a => 278, b => 310, p => false), (a => 5, b => 9, p => false), (a => 93, b => 97, p => false), (a => 181, b => 185, p => false), (a => 269, b => 273, p => false), (a => 13, b => 45, p => false), (a => 101, b => 133, p => false), (a => 189, b => 221, p => false), (a => 277, b => 309, p => false), (a => 7, b => 11, p => false), (a => 95, b => 99, p => false), (a => 183, b => 187, p => false), (a => 271, b => 275, p => false), (a => 15, b => 47, p => false), (a => 103, b => 135, p => false), (a => 191, b => 223, p => false), (a => 279, b => 311, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 16, b => 347, p => true), (a => 17, b => 346, p => true), (a => 18, b => 345, p => true), (a => 19, b => 344, p => true), (a => 20, b => 343, p => true), (a => 21, b => 342, p => true), (a => 22, b => 341, p => true), (a => 23, b => 340, p => true), (a => 24, b => 339, p => true), (a => 25, b => 338, p => true), (a => 26, b => 337, p => true), (a => 27, b => 336, p => true), (a => 28, b => 335, p => true), (a => 29, b => 334, p => true), (a => 30, b => 333, p => true), (a => 31, b => 332, p => true), (a => 32, b => 331, p => true), (a => 33, b => 330, p => true), (a => 34, b => 329, p => true), (a => 35, b => 328, p => true), (a => 36, b => 327, p => true), (a => 37, b => 326, p => true), (a => 38, b => 325, p => true), (a => 39, b => 324, p => true), (a => 40, b => 323, p => true), (a => 41, b => 322, p => true), (a => 42, b => 321, p => true), (a => 43, b => 320, p => true), (a => 48, b => 319, p => true), (a => 49, b => 318, p => true), (a => 50, b => 317, p => true), (a => 51, b => 316, p => true), (a => 52, b => 315, p => true), (a => 53, b => 314, p => true), (a => 54, b => 313, p => true), (a => 55, b => 312, p => true), (a => 56, b => 307, p => true), (a => 57, b => 306, p => true), (a => 58, b => 305, p => true), (a => 59, b => 304, p => true), (a => 60, b => 303, p => true), (a => 61, b => 302, p => true), (a => 62, b => 301, p => true), (a => 63, b => 300, p => true), (a => 64, b => 299, p => true), (a => 65, b => 298, p => true), (a => 66, b => 297, p => true), (a => 67, b => 296, p => true), (a => 68, b => 295, p => true), (a => 69, b => 294, p => true), (a => 70, b => 293, p => true), (a => 71, b => 292, p => true), (a => 72, b => 291, p => true), (a => 73, b => 290, p => true), (a => 74, b => 289, p => true), (a => 75, b => 288, p => true), (a => 76, b => 287, p => true), (a => 77, b => 286, p => true), (a => 78, b => 285, p => true), (a => 79, b => 284, p => true), (a => 80, b => 283, p => true), (a => 81, b => 282, p => true), (a => 82, b => 281, p => true), (a => 83, b => 280, p => true), (a => 84, b => 267, p => true), (a => 85, b => 266, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 90, b => 261, p => true), (a => 91, b => 260, p => true), (a => 104, b => 259, p => true), (a => 105, b => 258, p => true), (a => 106, b => 257, p => true), (a => 107, b => 256, p => true), (a => 108, b => 255, p => true), (a => 109, b => 254, p => true), (a => 110, b => 253, p => true), (a => 111, b => 252, p => true), (a => 112, b => 251, p => true), (a => 113, b => 250, p => true), (a => 114, b => 249, p => true), (a => 115, b => 248, p => true), (a => 116, b => 247, p => true), (a => 117, b => 246, p => true), (a => 118, b => 245, p => true), (a => 119, b => 244, p => true), (a => 120, b => 243, p => true), (a => 121, b => 242, p => true), (a => 122, b => 241, p => true), (a => 123, b => 240, p => true), (a => 124, b => 239, p => true), (a => 125, b => 238, p => true), (a => 126, b => 237, p => true), (a => 127, b => 236, p => true), (a => 128, b => 235, p => true), (a => 129, b => 234, p => true), (a => 130, b => 233, p => true), (a => 131, b => 232, p => true), (a => 136, b => 231, p => true), (a => 137, b => 230, p => true), (a => 138, b => 229, p => true), (a => 139, b => 228, p => true), (a => 140, b => 227, p => true), (a => 141, b => 226, p => true), (a => 142, b => 225, p => true), (a => 143, b => 224, p => true), (a => 144, b => 219, p => true), (a => 145, b => 218, p => true), (a => 146, b => 217, p => true), (a => 147, b => 216, p => true), (a => 148, b => 215, p => true), (a => 149, b => 214, p => true), (a => 150, b => 213, p => true), (a => 151, b => 212, p => true), (a => 152, b => 211, p => true), (a => 153, b => 210, p => true), (a => 154, b => 209, p => true), (a => 155, b => 208, p => true), (a => 156, b => 207, p => true), (a => 157, b => 206, p => true), (a => 158, b => 205, p => true), (a => 159, b => 204, p => true), (a => 160, b => 203, p => true), (a => 161, b => 202, p => true), (a => 162, b => 201, p => true), (a => 163, b => 200, p => true), (a => 164, b => 199, p => true), (a => 165, b => 198, p => true), (a => 166, b => 197, p => true), (a => 167, b => 196, p => true), (a => 168, b => 195, p => true), (a => 169, b => 194, p => true), (a => 170, b => 193, p => true), (a => 171, b => 192, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 2, b => 4, p => false), (a => 90, b => 92, p => false), (a => 178, b => 180, p => false), (a => 266, b => 268, p => false), (a => 6, b => 8, p => false), (a => 94, b => 96, p => false), (a => 182, b => 184, p => false), (a => 270, b => 272, p => false), (a => 10, b => 12, p => false), (a => 98, b => 100, p => false), (a => 186, b => 188, p => false), (a => 274, b => 276, p => false), (a => 14, b => 44, p => false), (a => 102, b => 132, p => false), (a => 190, b => 220, p => false), (a => 278, b => 308, p => false), (a => 3, b => 5, p => false), (a => 91, b => 93, p => false), (a => 179, b => 181, p => false), (a => 267, b => 269, p => false), (a => 7, b => 9, p => false), (a => 95, b => 97, p => false), (a => 183, b => 185, p => false), (a => 271, b => 273, p => false), (a => 11, b => 13, p => false), (a => 99, b => 101, p => false), (a => 187, b => 189, p => false), (a => 275, b => 277, p => false), (a => 15, b => 45, p => false), (a => 103, b => 133, p => false), (a => 191, b => 221, p => false), (a => 279, b => 309, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 16, b => 349, p => true), (a => 17, b => 348, p => true), (a => 18, b => 347, p => true), (a => 19, b => 346, p => true), (a => 20, b => 345, p => true), (a => 21, b => 344, p => true), (a => 22, b => 343, p => true), (a => 23, b => 342, p => true), (a => 24, b => 341, p => true), (a => 25, b => 340, p => true), (a => 26, b => 339, p => true), (a => 27, b => 338, p => true), (a => 28, b => 337, p => true), (a => 29, b => 336, p => true), (a => 30, b => 335, p => true), (a => 31, b => 334, p => true), (a => 32, b => 333, p => true), (a => 33, b => 332, p => true), (a => 34, b => 331, p => true), (a => 35, b => 330, p => true), (a => 36, b => 329, p => true), (a => 37, b => 328, p => true), (a => 38, b => 327, p => true), (a => 39, b => 326, p => true), (a => 40, b => 325, p => true), (a => 41, b => 324, p => true), (a => 42, b => 323, p => true), (a => 43, b => 322, p => true), (a => 46, b => 321, p => true), (a => 47, b => 320, p => true), (a => 48, b => 319, p => true), (a => 49, b => 318, p => true), (a => 50, b => 317, p => true), (a => 51, b => 316, p => true), (a => 52, b => 315, p => true), (a => 53, b => 314, p => true), (a => 54, b => 313, p => true), (a => 55, b => 312, p => true), (a => 56, b => 311, p => true), (a => 57, b => 310, p => true), (a => 58, b => 307, p => true), (a => 59, b => 306, p => true), (a => 60, b => 305, p => true), (a => 61, b => 304, p => true), (a => 62, b => 303, p => true), (a => 63, b => 302, p => true), (a => 64, b => 301, p => true), (a => 65, b => 300, p => true), (a => 66, b => 299, p => true), (a => 67, b => 298, p => true), (a => 68, b => 297, p => true), (a => 69, b => 296, p => true), (a => 70, b => 295, p => true), (a => 71, b => 294, p => true), (a => 72, b => 293, p => true), (a => 73, b => 292, p => true), (a => 74, b => 291, p => true), (a => 75, b => 290, p => true), (a => 76, b => 289, p => true), (a => 77, b => 288, p => true), (a => 78, b => 287, p => true), (a => 79, b => 286, p => true), (a => 80, b => 285, p => true), (a => 81, b => 284, p => true), (a => 82, b => 283, p => true), (a => 83, b => 282, p => true), (a => 84, b => 281, p => true), (a => 85, b => 280, p => true), (a => 86, b => 265, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 89, b => 262, p => true), (a => 104, b => 261, p => true), (a => 105, b => 260, p => true), (a => 106, b => 259, p => true), (a => 107, b => 258, p => true), (a => 108, b => 257, p => true), (a => 109, b => 256, p => true), (a => 110, b => 255, p => true), (a => 111, b => 254, p => true), (a => 112, b => 253, p => true), (a => 113, b => 252, p => true), (a => 114, b => 251, p => true), (a => 115, b => 250, p => true), (a => 116, b => 249, p => true), (a => 117, b => 248, p => true), (a => 118, b => 247, p => true), (a => 119, b => 246, p => true), (a => 120, b => 245, p => true), (a => 121, b => 244, p => true), (a => 122, b => 243, p => true), (a => 123, b => 242, p => true), (a => 124, b => 241, p => true), (a => 125, b => 240, p => true), (a => 126, b => 239, p => true), (a => 127, b => 238, p => true), (a => 128, b => 237, p => true), (a => 129, b => 236, p => true), (a => 130, b => 235, p => true), (a => 131, b => 234, p => true), (a => 134, b => 233, p => true), (a => 135, b => 232, p => true), (a => 136, b => 231, p => true), (a => 137, b => 230, p => true), (a => 138, b => 229, p => true), (a => 139, b => 228, p => true), (a => 140, b => 227, p => true), (a => 141, b => 226, p => true), (a => 142, b => 225, p => true), (a => 143, b => 224, p => true), (a => 144, b => 223, p => true), (a => 145, b => 222, p => true), (a => 146, b => 219, p => true), (a => 147, b => 218, p => true), (a => 148, b => 217, p => true), (a => 149, b => 216, p => true), (a => 150, b => 215, p => true), (a => 151, b => 214, p => true), (a => 152, b => 213, p => true), (a => 153, b => 212, p => true), (a => 154, b => 211, p => true), (a => 155, b => 210, p => true), (a => 156, b => 209, p => true), (a => 157, b => 208, p => true), (a => 158, b => 207, p => true), (a => 159, b => 206, p => true), (a => 160, b => 205, p => true), (a => 161, b => 204, p => true), (a => 162, b => 203, p => true), (a => 163, b => 202, p => true), (a => 164, b => 201, p => true), (a => 165, b => 200, p => true), (a => 166, b => 199, p => true), (a => 167, b => 198, p => true), (a => 168, b => 197, p => true), (a => 169, b => 196, p => true), (a => 170, b => 195, p => true), (a => 171, b => 194, p => true), (a => 172, b => 193, p => true), (a => 173, b => 192, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 1, b => 2, p => false), (a => 89, b => 90, p => false), (a => 177, b => 178, p => false), (a => 265, b => 266, p => false), (a => 3, b => 4, p => false), (a => 91, b => 92, p => false), (a => 179, b => 180, p => false), (a => 267, b => 268, p => false), (a => 5, b => 6, p => false), (a => 93, b => 94, p => false), (a => 181, b => 182, p => false), (a => 269, b => 270, p => false), (a => 7, b => 8, p => false), (a => 95, b => 96, p => false), (a => 183, b => 184, p => false), (a => 271, b => 272, p => false), (a => 9, b => 10, p => false), (a => 97, b => 98, p => false), (a => 185, b => 186, p => false), (a => 273, b => 274, p => false), (a => 11, b => 12, p => false), (a => 99, b => 100, p => false), (a => 187, b => 188, p => false), (a => 275, b => 276, p => false), (a => 13, b => 14, p => false), (a => 101, b => 102, p => false), (a => 189, b => 190, p => false), (a => 277, b => 278, p => false), (a => 15, b => 44, p => false), (a => 103, b => 132, p => false), (a => 191, b => 220, p => false), (a => 279, b => 308, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 22, b => 344, p => true), (a => 23, b => 343, p => true), (a => 24, b => 342, p => true), (a => 25, b => 341, p => true), (a => 26, b => 340, p => true), (a => 27, b => 339, p => true), (a => 28, b => 338, p => true), (a => 29, b => 337, p => true), (a => 30, b => 336, p => true), (a => 31, b => 335, p => true), (a => 32, b => 334, p => true), (a => 33, b => 333, p => true), (a => 34, b => 332, p => true), (a => 35, b => 331, p => true), (a => 36, b => 330, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 323, p => true), (a => 45, b => 322, p => true), (a => 46, b => 321, p => true), (a => 47, b => 320, p => true), (a => 48, b => 319, p => true), (a => 49, b => 318, p => true), (a => 50, b => 317, p => true), (a => 51, b => 316, p => true), (a => 52, b => 315, p => true), (a => 53, b => 314, p => true), (a => 54, b => 313, p => true), (a => 55, b => 312, p => true), (a => 56, b => 311, p => true), (a => 57, b => 310, p => true), (a => 58, b => 309, p => true), (a => 59, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 66, b => 300, p => true), (a => 67, b => 299, p => true), (a => 68, b => 298, p => true), (a => 69, b => 297, p => true), (a => 70, b => 296, p => true), (a => 71, b => 295, p => true), (a => 72, b => 294, p => true), (a => 73, b => 293, p => true), (a => 74, b => 292, p => true), (a => 75, b => 291, p => true), (a => 76, b => 290, p => true), (a => 77, b => 289, p => true), (a => 78, b => 288, p => true), (a => 79, b => 287, p => true), (a => 80, b => 286, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 110, b => 256, p => true), (a => 111, b => 255, p => true), (a => 112, b => 254, p => true), (a => 113, b => 253, p => true), (a => 114, b => 252, p => true), (a => 115, b => 251, p => true), (a => 116, b => 250, p => true), (a => 117, b => 249, p => true), (a => 118, b => 248, p => true), (a => 119, b => 247, p => true), (a => 120, b => 246, p => true), (a => 121, b => 245, p => true), (a => 122, b => 244, p => true), (a => 123, b => 243, p => true), (a => 124, b => 242, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 235, p => true), (a => 133, b => 234, p => true), (a => 134, b => 233, p => true), (a => 135, b => 232, p => true), (a => 136, b => 231, p => true), (a => 137, b => 230, p => true), (a => 138, b => 229, p => true), (a => 139, b => 228, p => true), (a => 140, b => 227, p => true), (a => 141, b => 226, p => true), (a => 142, b => 225, p => true), (a => 143, b => 224, p => true), (a => 144, b => 223, p => true), (a => 145, b => 222, p => true), (a => 146, b => 221, p => true), (a => 147, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 154, b => 212, p => true), (a => 155, b => 211, p => true), (a => 156, b => 210, p => true), (a => 157, b => 209, p => true), (a => 158, b => 208, p => true), (a => 159, b => 207, p => true), (a => 160, b => 206, p => true), (a => 161, b => 205, p => true), (a => 162, b => 204, p => true), (a => 163, b => 203, p => true), (a => 164, b => 202, p => true), (a => 165, b => 201, p => true), (a => 166, b => 200, p => true), (a => 167, b => 199, p => true), (a => 168, b => 198, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 96, p => false), (a => 184, b => 272, p => false), (a => 4, b => 92, p => false), (a => 180, b => 268, p => false), (a => 12, b => 100, p => false), (a => 188, b => 276, p => false), (a => 2, b => 90, p => false), (a => 178, b => 266, p => false), (a => 10, b => 98, p => false), (a => 186, b => 274, p => false), (a => 6, b => 94, p => false), (a => 182, b => 270, p => false), (a => 14, b => 102, p => false), (a => 190, b => 278, p => false), (a => 1, b => 89, p => false), (a => 177, b => 265, p => false), (a => 9, b => 97, p => false), (a => 185, b => 273, p => false), (a => 5, b => 93, p => false), (a => 181, b => 269, p => false), (a => 13, b => 101, p => false), (a => 189, b => 277, p => false), (a => 3, b => 91, p => false), (a => 179, b => 267, p => false), (a => 11, b => 99, p => false), (a => 187, b => 275, p => false), (a => 7, b => 95, p => false), (a => 183, b => 271, p => false), (a => 15, b => 103, p => false), (a => 191, b => 279, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 22, b => 344, p => true), (a => 23, b => 343, p => true), (a => 24, b => 342, p => true), (a => 25, b => 341, p => true), (a => 26, b => 340, p => true), (a => 27, b => 339, p => true), (a => 28, b => 338, p => true), (a => 29, b => 337, p => true), (a => 30, b => 336, p => true), (a => 31, b => 335, p => true), (a => 32, b => 334, p => true), (a => 33, b => 333, p => true), (a => 34, b => 332, p => true), (a => 35, b => 331, p => true), (a => 36, b => 330, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 323, p => true), (a => 44, b => 322, p => true), (a => 45, b => 321, p => true), (a => 46, b => 320, p => true), (a => 47, b => 319, p => true), (a => 48, b => 318, p => true), (a => 49, b => 317, p => true), (a => 50, b => 316, p => true), (a => 51, b => 315, p => true), (a => 52, b => 314, p => true), (a => 53, b => 313, p => true), (a => 54, b => 312, p => true), (a => 55, b => 311, p => true), (a => 56, b => 310, p => true), (a => 57, b => 309, p => true), (a => 58, b => 308, p => true), (a => 59, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 66, b => 300, p => true), (a => 67, b => 299, p => true), (a => 68, b => 298, p => true), (a => 69, b => 297, p => true), (a => 70, b => 296, p => true), (a => 71, b => 295, p => true), (a => 72, b => 294, p => true), (a => 73, b => 293, p => true), (a => 74, b => 292, p => true), (a => 75, b => 291, p => true), (a => 76, b => 290, p => true), (a => 77, b => 289, p => true), (a => 78, b => 288, p => true), (a => 79, b => 287, p => true), (a => 80, b => 286, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 264, p => true), (a => 88, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 110, b => 256, p => true), (a => 111, b => 255, p => true), (a => 112, b => 254, p => true), (a => 113, b => 253, p => true), (a => 114, b => 252, p => true), (a => 115, b => 251, p => true), (a => 116, b => 250, p => true), (a => 117, b => 249, p => true), (a => 118, b => 248, p => true), (a => 119, b => 247, p => true), (a => 120, b => 246, p => true), (a => 121, b => 245, p => true), (a => 122, b => 244, p => true), (a => 123, b => 243, p => true), (a => 124, b => 242, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 235, p => true), (a => 132, b => 234, p => true), (a => 133, b => 233, p => true), (a => 134, b => 232, p => true), (a => 135, b => 231, p => true), (a => 136, b => 230, p => true), (a => 137, b => 229, p => true), (a => 138, b => 228, p => true), (a => 139, b => 227, p => true), (a => 140, b => 226, p => true), (a => 141, b => 225, p => true), (a => 142, b => 224, p => true), (a => 143, b => 223, p => true), (a => 144, b => 222, p => true), (a => 145, b => 221, p => true), (a => 146, b => 220, p => true), (a => 147, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 154, b => 212, p => true), (a => 155, b => 211, p => true), (a => 156, b => 210, p => true), (a => 157, b => 209, p => true), (a => 158, b => 208, p => true), (a => 159, b => 207, p => true), (a => 160, b => 206, p => true), (a => 161, b => 205, p => true), (a => 162, b => 204, p => true), (a => 163, b => 203, p => true), (a => 164, b => 202, p => true), (a => 165, b => 201, p => true), (a => 166, b => 200, p => true), (a => 167, b => 199, p => true), (a => 168, b => 198, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 88, p => false), (a => 184, b => 264, p => false), (a => 12, b => 92, p => false), (a => 188, b => 268, p => false), (a => 10, b => 90, p => false), (a => 186, b => 266, p => false), (a => 14, b => 94, p => false), (a => 190, b => 270, p => false), (a => 9, b => 89, p => false), (a => 185, b => 265, p => false), (a => 13, b => 93, p => false), (a => 189, b => 269, p => false), (a => 11, b => 91, p => false), (a => 187, b => 267, p => false), (a => 15, b => 95, p => false), (a => 191, b => 271, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 4, b => 347, p => true), (a => 5, b => 346, p => true), (a => 6, b => 345, p => true), (a => 7, b => 344, p => true), (a => 16, b => 343, p => true), (a => 17, b => 342, p => true), (a => 18, b => 341, p => true), (a => 19, b => 340, p => true), (a => 20, b => 339, p => true), (a => 21, b => 338, p => true), (a => 22, b => 337, p => true), (a => 23, b => 336, p => true), (a => 24, b => 335, p => true), (a => 25, b => 334, p => true), (a => 26, b => 333, p => true), (a => 27, b => 332, p => true), (a => 28, b => 331, p => true), (a => 29, b => 330, p => true), (a => 30, b => 329, p => true), (a => 31, b => 328, p => true), (a => 32, b => 327, p => true), (a => 33, b => 326, p => true), (a => 34, b => 325, p => true), (a => 35, b => 324, p => true), (a => 36, b => 323, p => true), (a => 37, b => 322, p => true), (a => 38, b => 321, p => true), (a => 39, b => 320, p => true), (a => 40, b => 319, p => true), (a => 41, b => 318, p => true), (a => 42, b => 317, p => true), (a => 43, b => 316, p => true), (a => 44, b => 315, p => true), (a => 45, b => 314, p => true), (a => 46, b => 313, p => true), (a => 47, b => 312, p => true), (a => 48, b => 311, p => true), (a => 49, b => 310, p => true), (a => 50, b => 309, p => true), (a => 51, b => 308, p => true), (a => 52, b => 307, p => true), (a => 53, b => 306, p => true), (a => 54, b => 305, p => true), (a => 55, b => 304, p => true), (a => 56, b => 303, p => true), (a => 57, b => 302, p => true), (a => 58, b => 301, p => true), (a => 59, b => 300, p => true), (a => 60, b => 299, p => true), (a => 61, b => 298, p => true), (a => 62, b => 297, p => true), (a => 63, b => 296, p => true), (a => 64, b => 295, p => true), (a => 65, b => 294, p => true), (a => 66, b => 293, p => true), (a => 67, b => 292, p => true), (a => 68, b => 291, p => true), (a => 69, b => 290, p => true), (a => 70, b => 289, p => true), (a => 71, b => 288, p => true), (a => 72, b => 287, p => true), (a => 73, b => 286, p => true), (a => 74, b => 285, p => true), (a => 75, b => 284, p => true), (a => 76, b => 283, p => true), (a => 77, b => 282, p => true), (a => 78, b => 281, p => true), (a => 79, b => 280, p => true), (a => 80, b => 279, p => true), (a => 81, b => 278, p => true), (a => 82, b => 277, p => true), (a => 83, b => 276, p => true), (a => 84, b => 275, p => true), (a => 85, b => 274, p => true), (a => 86, b => 273, p => true), (a => 87, b => 272, p => true), (a => 96, b => 263, p => true), (a => 97, b => 262, p => true), (a => 98, b => 261, p => true), (a => 99, b => 260, p => true), (a => 100, b => 259, p => true), (a => 101, b => 258, p => true), (a => 102, b => 257, p => true), (a => 103, b => 256, p => true), (a => 104, b => 255, p => true), (a => 105, b => 254, p => true), (a => 106, b => 253, p => true), (a => 107, b => 252, p => true), (a => 108, b => 251, p => true), (a => 109, b => 250, p => true), (a => 110, b => 249, p => true), (a => 111, b => 248, p => true), (a => 112, b => 247, p => true), (a => 113, b => 246, p => true), (a => 114, b => 245, p => true), (a => 115, b => 244, p => true), (a => 116, b => 243, p => true), (a => 117, b => 242, p => true), (a => 118, b => 241, p => true), (a => 119, b => 240, p => true), (a => 120, b => 239, p => true), (a => 121, b => 238, p => true), (a => 122, b => 237, p => true), (a => 123, b => 236, p => true), (a => 124, b => 235, p => true), (a => 125, b => 234, p => true), (a => 126, b => 233, p => true), (a => 127, b => 232, p => true), (a => 128, b => 231, p => true), (a => 129, b => 230, p => true), (a => 130, b => 229, p => true), (a => 131, b => 228, p => true), (a => 132, b => 227, p => true), (a => 133, b => 226, p => true), (a => 134, b => 225, p => true), (a => 135, b => 224, p => true), (a => 136, b => 223, p => true), (a => 137, b => 222, p => true), (a => 138, b => 221, p => true), (a => 139, b => 220, p => true), (a => 140, b => 219, p => true), (a => 141, b => 218, p => true), (a => 142, b => 217, p => true), (a => 143, b => 216, p => true), (a => 144, b => 215, p => true), (a => 145, b => 214, p => true), (a => 146, b => 213, p => true), (a => 147, b => 212, p => true), (a => 148, b => 211, p => true), (a => 149, b => 210, p => true), (a => 150, b => 209, p => true), (a => 151, b => 208, p => true), (a => 152, b => 207, p => true), (a => 153, b => 206, p => true), (a => 154, b => 205, p => true), (a => 155, b => 204, p => true), (a => 156, b => 203, p => true), (a => 157, b => 202, p => true), (a => 158, b => 201, p => true), (a => 159, b => 200, p => true), (a => 160, b => 199, p => true), (a => 161, b => 198, p => true), (a => 162, b => 197, p => true), (a => 163, b => 196, p => true), (a => 164, b => 195, p => true), (a => 165, b => 194, p => true), (a => 166, b => 193, p => true), (a => 167, b => 192, p => true), (a => 168, b => 183, p => true), (a => 169, b => 182, p => true), (a => 170, b => 181, p => true), (a => 171, b => 180, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 4, b => 8, p => false), (a => 180, b => 184, p => false), (a => 12, b => 88, p => false), (a => 188, b => 264, p => false), (a => 6, b => 10, p => false), (a => 182, b => 186, p => false), (a => 14, b => 90, p => false), (a => 190, b => 266, p => false), (a => 5, b => 9, p => false), (a => 181, b => 185, p => false), (a => 13, b => 89, p => false), (a => 189, b => 265, p => false), (a => 7, b => 11, p => false), (a => 183, b => 187, p => false), (a => 15, b => 91, p => false), (a => 191, b => 267, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 16, b => 347, p => true), (a => 17, b => 346, p => true), (a => 18, b => 345, p => true), (a => 19, b => 344, p => true), (a => 20, b => 343, p => true), (a => 21, b => 342, p => true), (a => 22, b => 341, p => true), (a => 23, b => 340, p => true), (a => 24, b => 339, p => true), (a => 25, b => 338, p => true), (a => 26, b => 337, p => true), (a => 27, b => 336, p => true), (a => 28, b => 335, p => true), (a => 29, b => 334, p => true), (a => 30, b => 333, p => true), (a => 31, b => 332, p => true), (a => 32, b => 331, p => true), (a => 33, b => 330, p => true), (a => 34, b => 329, p => true), (a => 35, b => 328, p => true), (a => 36, b => 327, p => true), (a => 37, b => 326, p => true), (a => 38, b => 325, p => true), (a => 39, b => 324, p => true), (a => 40, b => 323, p => true), (a => 41, b => 322, p => true), (a => 42, b => 321, p => true), (a => 43, b => 320, p => true), (a => 44, b => 319, p => true), (a => 45, b => 318, p => true), (a => 46, b => 317, p => true), (a => 47, b => 316, p => true), (a => 48, b => 315, p => true), (a => 49, b => 314, p => true), (a => 50, b => 313, p => true), (a => 51, b => 312, p => true), (a => 52, b => 311, p => true), (a => 53, b => 310, p => true), (a => 54, b => 309, p => true), (a => 55, b => 308, p => true), (a => 56, b => 307, p => true), (a => 57, b => 306, p => true), (a => 58, b => 305, p => true), (a => 59, b => 304, p => true), (a => 60, b => 303, p => true), (a => 61, b => 302, p => true), (a => 62, b => 301, p => true), (a => 63, b => 300, p => true), (a => 64, b => 299, p => true), (a => 65, b => 298, p => true), (a => 66, b => 297, p => true), (a => 67, b => 296, p => true), (a => 68, b => 295, p => true), (a => 69, b => 294, p => true), (a => 70, b => 293, p => true), (a => 71, b => 292, p => true), (a => 72, b => 291, p => true), (a => 73, b => 290, p => true), (a => 74, b => 289, p => true), (a => 75, b => 288, p => true), (a => 76, b => 287, p => true), (a => 77, b => 286, p => true), (a => 78, b => 285, p => true), (a => 79, b => 284, p => true), (a => 80, b => 283, p => true), (a => 81, b => 282, p => true), (a => 82, b => 281, p => true), (a => 83, b => 280, p => true), (a => 84, b => 279, p => true), (a => 85, b => 278, p => true), (a => 86, b => 277, p => true), (a => 87, b => 276, p => true), (a => 92, b => 275, p => true), (a => 93, b => 274, p => true), (a => 94, b => 273, p => true), (a => 95, b => 272, p => true), (a => 96, b => 271, p => true), (a => 97, b => 270, p => true), (a => 98, b => 269, p => true), (a => 99, b => 268, p => true), (a => 100, b => 263, p => true), (a => 101, b => 262, p => true), (a => 102, b => 261, p => true), (a => 103, b => 260, p => true), (a => 104, b => 259, p => true), (a => 105, b => 258, p => true), (a => 106, b => 257, p => true), (a => 107, b => 256, p => true), (a => 108, b => 255, p => true), (a => 109, b => 254, p => true), (a => 110, b => 253, p => true), (a => 111, b => 252, p => true), (a => 112, b => 251, p => true), (a => 113, b => 250, p => true), (a => 114, b => 249, p => true), (a => 115, b => 248, p => true), (a => 116, b => 247, p => true), (a => 117, b => 246, p => true), (a => 118, b => 245, p => true), (a => 119, b => 244, p => true), (a => 120, b => 243, p => true), (a => 121, b => 242, p => true), (a => 122, b => 241, p => true), (a => 123, b => 240, p => true), (a => 124, b => 239, p => true), (a => 125, b => 238, p => true), (a => 126, b => 237, p => true), (a => 127, b => 236, p => true), (a => 128, b => 235, p => true), (a => 129, b => 234, p => true), (a => 130, b => 233, p => true), (a => 131, b => 232, p => true), (a => 132, b => 231, p => true), (a => 133, b => 230, p => true), (a => 134, b => 229, p => true), (a => 135, b => 228, p => true), (a => 136, b => 227, p => true), (a => 137, b => 226, p => true), (a => 138, b => 225, p => true), (a => 139, b => 224, p => true), (a => 140, b => 223, p => true), (a => 141, b => 222, p => true), (a => 142, b => 221, p => true), (a => 143, b => 220, p => true), (a => 144, b => 219, p => true), (a => 145, b => 218, p => true), (a => 146, b => 217, p => true), (a => 147, b => 216, p => true), (a => 148, b => 215, p => true), (a => 149, b => 214, p => true), (a => 150, b => 213, p => true), (a => 151, b => 212, p => true), (a => 152, b => 211, p => true), (a => 153, b => 210, p => true), (a => 154, b => 209, p => true), (a => 155, b => 208, p => true), (a => 156, b => 207, p => true), (a => 157, b => 206, p => true), (a => 158, b => 205, p => true), (a => 159, b => 204, p => true), (a => 160, b => 203, p => true), (a => 161, b => 202, p => true), (a => 162, b => 201, p => true), (a => 163, b => 200, p => true), (a => 164, b => 199, p => true), (a => 165, b => 198, p => true), (a => 166, b => 197, p => true), (a => 167, b => 196, p => true), (a => 168, b => 195, p => true), (a => 169, b => 194, p => true), (a => 170, b => 193, p => true), (a => 171, b => 192, p => true), (a => 172, b => 179, p => true), (a => 173, b => 178, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 2, b => 4, p => false), (a => 178, b => 180, p => false), (a => 6, b => 8, p => false), (a => 182, b => 184, p => false), (a => 10, b => 12, p => false), (a => 186, b => 188, p => false), (a => 14, b => 88, p => false), (a => 190, b => 264, p => false), (a => 3, b => 5, p => false), (a => 179, b => 181, p => false), (a => 7, b => 9, p => false), (a => 183, b => 185, p => false), (a => 11, b => 13, p => false), (a => 187, b => 189, p => false), (a => 15, b => 89, p => false), (a => 191, b => 265, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 16, b => 349, p => true), (a => 17, b => 348, p => true), (a => 18, b => 347, p => true), (a => 19, b => 346, p => true), (a => 20, b => 345, p => true), (a => 21, b => 344, p => true), (a => 22, b => 343, p => true), (a => 23, b => 342, p => true), (a => 24, b => 341, p => true), (a => 25, b => 340, p => true), (a => 26, b => 339, p => true), (a => 27, b => 338, p => true), (a => 28, b => 337, p => true), (a => 29, b => 336, p => true), (a => 30, b => 335, p => true), (a => 31, b => 334, p => true), (a => 32, b => 333, p => true), (a => 33, b => 332, p => true), (a => 34, b => 331, p => true), (a => 35, b => 330, p => true), (a => 36, b => 329, p => true), (a => 37, b => 328, p => true), (a => 38, b => 327, p => true), (a => 39, b => 326, p => true), (a => 40, b => 325, p => true), (a => 41, b => 324, p => true), (a => 42, b => 323, p => true), (a => 43, b => 322, p => true), (a => 44, b => 321, p => true), (a => 45, b => 320, p => true), (a => 46, b => 319, p => true), (a => 47, b => 318, p => true), (a => 48, b => 317, p => true), (a => 49, b => 316, p => true), (a => 50, b => 315, p => true), (a => 51, b => 314, p => true), (a => 52, b => 313, p => true), (a => 53, b => 312, p => true), (a => 54, b => 311, p => true), (a => 55, b => 310, p => true), (a => 56, b => 309, p => true), (a => 57, b => 308, p => true), (a => 58, b => 307, p => true), (a => 59, b => 306, p => true), (a => 60, b => 305, p => true), (a => 61, b => 304, p => true), (a => 62, b => 303, p => true), (a => 63, b => 302, p => true), (a => 64, b => 301, p => true), (a => 65, b => 300, p => true), (a => 66, b => 299, p => true), (a => 67, b => 298, p => true), (a => 68, b => 297, p => true), (a => 69, b => 296, p => true), (a => 70, b => 295, p => true), (a => 71, b => 294, p => true), (a => 72, b => 293, p => true), (a => 73, b => 292, p => true), (a => 74, b => 291, p => true), (a => 75, b => 290, p => true), (a => 76, b => 289, p => true), (a => 77, b => 288, p => true), (a => 78, b => 287, p => true), (a => 79, b => 286, p => true), (a => 80, b => 285, p => true), (a => 81, b => 284, p => true), (a => 82, b => 283, p => true), (a => 83, b => 282, p => true), (a => 84, b => 281, p => true), (a => 85, b => 280, p => true), (a => 86, b => 279, p => true), (a => 87, b => 278, p => true), (a => 90, b => 277, p => true), (a => 91, b => 276, p => true), (a => 92, b => 275, p => true), (a => 93, b => 274, p => true), (a => 94, b => 273, p => true), (a => 95, b => 272, p => true), (a => 96, b => 271, p => true), (a => 97, b => 270, p => true), (a => 98, b => 269, p => true), (a => 99, b => 268, p => true), (a => 100, b => 267, p => true), (a => 101, b => 266, p => true), (a => 102, b => 263, p => true), (a => 103, b => 262, p => true), (a => 104, b => 261, p => true), (a => 105, b => 260, p => true), (a => 106, b => 259, p => true), (a => 107, b => 258, p => true), (a => 108, b => 257, p => true), (a => 109, b => 256, p => true), (a => 110, b => 255, p => true), (a => 111, b => 254, p => true), (a => 112, b => 253, p => true), (a => 113, b => 252, p => true), (a => 114, b => 251, p => true), (a => 115, b => 250, p => true), (a => 116, b => 249, p => true), (a => 117, b => 248, p => true), (a => 118, b => 247, p => true), (a => 119, b => 246, p => true), (a => 120, b => 245, p => true), (a => 121, b => 244, p => true), (a => 122, b => 243, p => true), (a => 123, b => 242, p => true), (a => 124, b => 241, p => true), (a => 125, b => 240, p => true), (a => 126, b => 239, p => true), (a => 127, b => 238, p => true), (a => 128, b => 237, p => true), (a => 129, b => 236, p => true), (a => 130, b => 235, p => true), (a => 131, b => 234, p => true), (a => 132, b => 233, p => true), (a => 133, b => 232, p => true), (a => 134, b => 231, p => true), (a => 135, b => 230, p => true), (a => 136, b => 229, p => true), (a => 137, b => 228, p => true), (a => 138, b => 227, p => true), (a => 139, b => 226, p => true), (a => 140, b => 225, p => true), (a => 141, b => 224, p => true), (a => 142, b => 223, p => true), (a => 143, b => 222, p => true), (a => 144, b => 221, p => true), (a => 145, b => 220, p => true), (a => 146, b => 219, p => true), (a => 147, b => 218, p => true), (a => 148, b => 217, p => true), (a => 149, b => 216, p => true), (a => 150, b => 215, p => true), (a => 151, b => 214, p => true), (a => 152, b => 213, p => true), (a => 153, b => 212, p => true), (a => 154, b => 211, p => true), (a => 155, b => 210, p => true), (a => 156, b => 209, p => true), (a => 157, b => 208, p => true), (a => 158, b => 207, p => true), (a => 159, b => 206, p => true), (a => 160, b => 205, p => true), (a => 161, b => 204, p => true), (a => 162, b => 203, p => true), (a => 163, b => 202, p => true), (a => 164, b => 201, p => true), (a => 165, b => 200, p => true), (a => 166, b => 199, p => true), (a => 167, b => 198, p => true), (a => 168, b => 197, p => true), (a => 169, b => 196, p => true), (a => 170, b => 195, p => true), (a => 171, b => 194, p => true), (a => 172, b => 193, p => true), (a => 173, b => 192, p => true), (a => 174, b => 177, p => true), (a => 175, b => 176, p => true)),
        ((a    => 1, b => 2, p => false), (a => 177, b => 178, p => false), (a => 3, b => 4, p => false), (a => 179, b => 180, p => false), (a => 5, b => 6, p => false), (a => 181, b => 182, p => false), (a => 7, b => 8, p => false), (a => 183, b => 184, p => false), (a => 9, b => 10, p => false), (a => 185, b => 186, p => false), (a => 11, b => 12, p => false), (a => 187, b => 188, p => false), (a => 13, b => 14, p => false), (a => 189, b => 190, p => false), (a => 15, b => 88, p => false), (a => 191, b => 264, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 22, b => 344, p => true), (a => 23, b => 343, p => true), (a => 24, b => 342, p => true), (a => 25, b => 341, p => true), (a => 26, b => 340, p => true), (a => 27, b => 339, p => true), (a => 28, b => 338, p => true), (a => 29, b => 337, p => true), (a => 30, b => 336, p => true), (a => 31, b => 335, p => true), (a => 32, b => 334, p => true), (a => 33, b => 333, p => true), (a => 34, b => 332, p => true), (a => 35, b => 331, p => true), (a => 36, b => 330, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 323, p => true), (a => 44, b => 322, p => true), (a => 45, b => 321, p => true), (a => 46, b => 320, p => true), (a => 47, b => 319, p => true), (a => 48, b => 318, p => true), (a => 49, b => 317, p => true), (a => 50, b => 316, p => true), (a => 51, b => 315, p => true), (a => 52, b => 314, p => true), (a => 53, b => 313, p => true), (a => 54, b => 312, p => true), (a => 55, b => 311, p => true), (a => 56, b => 310, p => true), (a => 57, b => 309, p => true), (a => 58, b => 308, p => true), (a => 59, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 66, b => 300, p => true), (a => 67, b => 299, p => true), (a => 68, b => 298, p => true), (a => 69, b => 297, p => true), (a => 70, b => 296, p => true), (a => 71, b => 295, p => true), (a => 72, b => 294, p => true), (a => 73, b => 293, p => true), (a => 74, b => 292, p => true), (a => 75, b => 291, p => true), (a => 76, b => 290, p => true), (a => 77, b => 289, p => true), (a => 78, b => 288, p => true), (a => 79, b => 287, p => true), (a => 80, b => 286, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 279, p => true), (a => 89, b => 278, p => true), (a => 90, b => 277, p => true), (a => 91, b => 276, p => true), (a => 92, b => 275, p => true), (a => 93, b => 274, p => true), (a => 94, b => 273, p => true), (a => 95, b => 272, p => true), (a => 96, b => 271, p => true), (a => 97, b => 270, p => true), (a => 98, b => 269, p => true), (a => 99, b => 268, p => true), (a => 100, b => 267, p => true), (a => 101, b => 266, p => true), (a => 102, b => 265, p => true), (a => 103, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 110, b => 256, p => true), (a => 111, b => 255, p => true), (a => 112, b => 254, p => true), (a => 113, b => 253, p => true), (a => 114, b => 252, p => true), (a => 115, b => 251, p => true), (a => 116, b => 250, p => true), (a => 117, b => 249, p => true), (a => 118, b => 248, p => true), (a => 119, b => 247, p => true), (a => 120, b => 246, p => true), (a => 121, b => 245, p => true), (a => 122, b => 244, p => true), (a => 123, b => 243, p => true), (a => 124, b => 242, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 235, p => true), (a => 132, b => 234, p => true), (a => 133, b => 233, p => true), (a => 134, b => 232, p => true), (a => 135, b => 231, p => true), (a => 136, b => 230, p => true), (a => 137, b => 229, p => true), (a => 138, b => 228, p => true), (a => 139, b => 227, p => true), (a => 140, b => 226, p => true), (a => 141, b => 225, p => true), (a => 142, b => 224, p => true), (a => 143, b => 223, p => true), (a => 144, b => 222, p => true), (a => 145, b => 221, p => true), (a => 146, b => 220, p => true), (a => 147, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 154, b => 212, p => true), (a => 155, b => 211, p => true), (a => 156, b => 210, p => true), (a => 157, b => 209, p => true), (a => 158, b => 208, p => true), (a => 159, b => 207, p => true), (a => 160, b => 206, p => true), (a => 161, b => 205, p => true), (a => 162, b => 204, p => true), (a => 163, b => 203, p => true), (a => 164, b => 202, p => true), (a => 165, b => 201, p => true), (a => 166, b => 200, p => true), (a => 167, b => 199, p => true), (a => 168, b => 198, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 184, p => false), (a => 4, b => 180, p => false), (a => 12, b => 188, p => false), (a => 2, b => 178, p => false), (a => 10, b => 186, p => false), (a => 6, b => 182, p => false), (a => 14, b => 190, p => false), (a => 1, b => 177, p => false), (a => 9, b => 185, p => false), (a => 5, b => 181, p => false), (a => 13, b => 189, p => false), (a => 3, b => 179, p => false), (a => 11, b => 187, p => false), (a => 7, b => 183, p => false), (a => 15, b => 191, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 22, b => 344, p => true), (a => 23, b => 343, p => true), (a => 24, b => 342, p => true), (a => 25, b => 341, p => true), (a => 26, b => 340, p => true), (a => 27, b => 339, p => true), (a => 28, b => 338, p => true), (a => 29, b => 337, p => true), (a => 30, b => 336, p => true), (a => 31, b => 335, p => true), (a => 32, b => 334, p => true), (a => 33, b => 333, p => true), (a => 34, b => 332, p => true), (a => 35, b => 331, p => true), (a => 36, b => 330, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 323, p => true), (a => 44, b => 322, p => true), (a => 45, b => 321, p => true), (a => 46, b => 320, p => true), (a => 47, b => 319, p => true), (a => 48, b => 318, p => true), (a => 49, b => 317, p => true), (a => 50, b => 316, p => true), (a => 51, b => 315, p => true), (a => 52, b => 314, p => true), (a => 53, b => 313, p => true), (a => 54, b => 312, p => true), (a => 55, b => 311, p => true), (a => 56, b => 310, p => true), (a => 57, b => 309, p => true), (a => 58, b => 308, p => true), (a => 59, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 66, b => 300, p => true), (a => 67, b => 299, p => true), (a => 68, b => 298, p => true), (a => 69, b => 297, p => true), (a => 70, b => 296, p => true), (a => 71, b => 295, p => true), (a => 72, b => 294, p => true), (a => 73, b => 293, p => true), (a => 74, b => 292, p => true), (a => 75, b => 291, p => true), (a => 76, b => 290, p => true), (a => 77, b => 289, p => true), (a => 78, b => 288, p => true), (a => 79, b => 287, p => true), (a => 80, b => 286, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 279, p => true), (a => 88, b => 278, p => true), (a => 89, b => 277, p => true), (a => 90, b => 276, p => true), (a => 91, b => 275, p => true), (a => 92, b => 274, p => true), (a => 93, b => 273, p => true), (a => 94, b => 272, p => true), (a => 95, b => 271, p => true), (a => 96, b => 270, p => true), (a => 97, b => 269, p => true), (a => 98, b => 268, p => true), (a => 99, b => 267, p => true), (a => 100, b => 266, p => true), (a => 101, b => 265, p => true), (a => 102, b => 264, p => true), (a => 103, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 110, b => 256, p => true), (a => 111, b => 255, p => true), (a => 112, b => 254, p => true), (a => 113, b => 253, p => true), (a => 114, b => 252, p => true), (a => 115, b => 251, p => true), (a => 116, b => 250, p => true), (a => 117, b => 249, p => true), (a => 118, b => 248, p => true), (a => 119, b => 247, p => true), (a => 120, b => 246, p => true), (a => 121, b => 245, p => true), (a => 122, b => 244, p => true), (a => 123, b => 243, p => true), (a => 124, b => 242, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 235, p => true), (a => 132, b => 234, p => true), (a => 133, b => 233, p => true), (a => 134, b => 232, p => true), (a => 135, b => 231, p => true), (a => 136, b => 230, p => true), (a => 137, b => 229, p => true), (a => 138, b => 228, p => true), (a => 139, b => 227, p => true), (a => 140, b => 226, p => true), (a => 141, b => 225, p => true), (a => 142, b => 224, p => true), (a => 143, b => 223, p => true), (a => 144, b => 222, p => true), (a => 145, b => 221, p => true), (a => 146, b => 220, p => true), (a => 147, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 154, b => 212, p => true), (a => 155, b => 211, p => true), (a => 156, b => 210, p => true), (a => 157, b => 209, p => true), (a => 158, b => 208, p => true), (a => 159, b => 207, p => true), (a => 160, b => 206, p => true), (a => 161, b => 205, p => true), (a => 162, b => 204, p => true), (a => 163, b => 203, p => true), (a => 164, b => 202, p => true), (a => 165, b => 201, p => true), (a => 166, b => 200, p => true), (a => 167, b => 199, p => true), (a => 168, b => 198, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 176, p => true)),
        ((a    => 8, b => 176, p => false), (a => 12, b => 180, p => false), (a => 10, b => 178, p => false), (a => 14, b => 182, p => false), (a => 9, b => 177, p => false), (a => 13, b => 181, p => false), (a => 11, b => 179, p => false), (a => 15, b => 183, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 4, b => 347, p => true), (a => 5, b => 346, p => true), (a => 6, b => 345, p => true), (a => 7, b => 344, p => true), (a => 16, b => 343, p => true), (a => 17, b => 342, p => true), (a => 18, b => 341, p => true), (a => 19, b => 340, p => true), (a => 20, b => 339, p => true), (a => 21, b => 338, p => true), (a => 22, b => 337, p => true), (a => 23, b => 336, p => true), (a => 24, b => 335, p => true), (a => 25, b => 334, p => true), (a => 26, b => 333, p => true), (a => 27, b => 332, p => true), (a => 28, b => 331, p => true), (a => 29, b => 330, p => true), (a => 30, b => 329, p => true), (a => 31, b => 328, p => true), (a => 32, b => 327, p => true), (a => 33, b => 326, p => true), (a => 34, b => 325, p => true), (a => 35, b => 324, p => true), (a => 36, b => 323, p => true), (a => 37, b => 322, p => true), (a => 38, b => 321, p => true), (a => 39, b => 320, p => true), (a => 40, b => 319, p => true), (a => 41, b => 318, p => true), (a => 42, b => 317, p => true), (a => 43, b => 316, p => true), (a => 44, b => 315, p => true), (a => 45, b => 314, p => true), (a => 46, b => 313, p => true), (a => 47, b => 312, p => true), (a => 48, b => 311, p => true), (a => 49, b => 310, p => true), (a => 50, b => 309, p => true), (a => 51, b => 308, p => true), (a => 52, b => 307, p => true), (a => 53, b => 306, p => true), (a => 54, b => 305, p => true), (a => 55, b => 304, p => true), (a => 56, b => 303, p => true), (a => 57, b => 302, p => true), (a => 58, b => 301, p => true), (a => 59, b => 300, p => true), (a => 60, b => 299, p => true), (a => 61, b => 298, p => true), (a => 62, b => 297, p => true), (a => 63, b => 296, p => true), (a => 64, b => 295, p => true), (a => 65, b => 294, p => true), (a => 66, b => 293, p => true), (a => 67, b => 292, p => true), (a => 68, b => 291, p => true), (a => 69, b => 290, p => true), (a => 70, b => 289, p => true), (a => 71, b => 288, p => true), (a => 72, b => 287, p => true), (a => 73, b => 286, p => true), (a => 74, b => 285, p => true), (a => 75, b => 284, p => true), (a => 76, b => 283, p => true), (a => 77, b => 282, p => true), (a => 78, b => 281, p => true), (a => 79, b => 280, p => true), (a => 80, b => 279, p => true), (a => 81, b => 278, p => true), (a => 82, b => 277, p => true), (a => 83, b => 276, p => true), (a => 84, b => 275, p => true), (a => 85, b => 274, p => true), (a => 86, b => 273, p => true), (a => 87, b => 272, p => true), (a => 88, b => 271, p => true), (a => 89, b => 270, p => true), (a => 90, b => 269, p => true), (a => 91, b => 268, p => true), (a => 92, b => 267, p => true), (a => 93, b => 266, p => true), (a => 94, b => 265, p => true), (a => 95, b => 264, p => true), (a => 96, b => 263, p => true), (a => 97, b => 262, p => true), (a => 98, b => 261, p => true), (a => 99, b => 260, p => true), (a => 100, b => 259, p => true), (a => 101, b => 258, p => true), (a => 102, b => 257, p => true), (a => 103, b => 256, p => true), (a => 104, b => 255, p => true), (a => 105, b => 254, p => true), (a => 106, b => 253, p => true), (a => 107, b => 252, p => true), (a => 108, b => 251, p => true), (a => 109, b => 250, p => true), (a => 110, b => 249, p => true), (a => 111, b => 248, p => true), (a => 112, b => 247, p => true), (a => 113, b => 246, p => true), (a => 114, b => 245, p => true), (a => 115, b => 244, p => true), (a => 116, b => 243, p => true), (a => 117, b => 242, p => true), (a => 118, b => 241, p => true), (a => 119, b => 240, p => true), (a => 120, b => 239, p => true), (a => 121, b => 238, p => true), (a => 122, b => 237, p => true), (a => 123, b => 236, p => true), (a => 124, b => 235, p => true), (a => 125, b => 234, p => true), (a => 126, b => 233, p => true), (a => 127, b => 232, p => true), (a => 128, b => 231, p => true), (a => 129, b => 230, p => true), (a => 130, b => 229, p => true), (a => 131, b => 228, p => true), (a => 132, b => 227, p => true), (a => 133, b => 226, p => true), (a => 134, b => 225, p => true), (a => 135, b => 224, p => true), (a => 136, b => 223, p => true), (a => 137, b => 222, p => true), (a => 138, b => 221, p => true), (a => 139, b => 220, p => true), (a => 140, b => 219, p => true), (a => 141, b => 218, p => true), (a => 142, b => 217, p => true), (a => 143, b => 216, p => true), (a => 144, b => 215, p => true), (a => 145, b => 214, p => true), (a => 146, b => 213, p => true), (a => 147, b => 212, p => true), (a => 148, b => 211, p => true), (a => 149, b => 210, p => true), (a => 150, b => 209, p => true), (a => 151, b => 208, p => true), (a => 152, b => 207, p => true), (a => 153, b => 206, p => true), (a => 154, b => 205, p => true), (a => 155, b => 204, p => true), (a => 156, b => 203, p => true), (a => 157, b => 202, p => true), (a => 158, b => 201, p => true), (a => 159, b => 200, p => true), (a => 160, b => 199, p => true), (a => 161, b => 198, p => true), (a => 162, b => 197, p => true), (a => 163, b => 196, p => true), (a => 164, b => 195, p => true), (a => 165, b => 194, p => true), (a => 166, b => 193, p => true), (a => 167, b => 192, p => true), (a => 168, b => 191, p => true), (a => 169, b => 190, p => true), (a => 170, b => 189, p => true), (a => 171, b => 188, p => true), (a => 172, b => 187, p => true), (a => 173, b => 186, p => true), (a => 174, b => 185, p => true), (a => 175, b => 184, p => true)),
        ((a    => 4, b => 8, p => false), (a => 12, b => 176, p => false), (a => 6, b => 10, p => false), (a => 14, b => 178, p => false), (a => 5, b => 9, p => false), (a => 13, b => 177, p => false), (a => 7, b => 11, p => false), (a => 15, b => 179, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 2, b => 349, p => true), (a => 3, b => 348, p => true), (a => 16, b => 347, p => true), (a => 17, b => 346, p => true), (a => 18, b => 345, p => true), (a => 19, b => 344, p => true), (a => 20, b => 343, p => true), (a => 21, b => 342, p => true), (a => 22, b => 341, p => true), (a => 23, b => 340, p => true), (a => 24, b => 339, p => true), (a => 25, b => 338, p => true), (a => 26, b => 337, p => true), (a => 27, b => 336, p => true), (a => 28, b => 335, p => true), (a => 29, b => 334, p => true), (a => 30, b => 333, p => true), (a => 31, b => 332, p => true), (a => 32, b => 331, p => true), (a => 33, b => 330, p => true), (a => 34, b => 329, p => true), (a => 35, b => 328, p => true), (a => 36, b => 327, p => true), (a => 37, b => 326, p => true), (a => 38, b => 325, p => true), (a => 39, b => 324, p => true), (a => 40, b => 323, p => true), (a => 41, b => 322, p => true), (a => 42, b => 321, p => true), (a => 43, b => 320, p => true), (a => 44, b => 319, p => true), (a => 45, b => 318, p => true), (a => 46, b => 317, p => true), (a => 47, b => 316, p => true), (a => 48, b => 315, p => true), (a => 49, b => 314, p => true), (a => 50, b => 313, p => true), (a => 51, b => 312, p => true), (a => 52, b => 311, p => true), (a => 53, b => 310, p => true), (a => 54, b => 309, p => true), (a => 55, b => 308, p => true), (a => 56, b => 307, p => true), (a => 57, b => 306, p => true), (a => 58, b => 305, p => true), (a => 59, b => 304, p => true), (a => 60, b => 303, p => true), (a => 61, b => 302, p => true), (a => 62, b => 301, p => true), (a => 63, b => 300, p => true), (a => 64, b => 299, p => true), (a => 65, b => 298, p => true), (a => 66, b => 297, p => true), (a => 67, b => 296, p => true), (a => 68, b => 295, p => true), (a => 69, b => 294, p => true), (a => 70, b => 293, p => true), (a => 71, b => 292, p => true), (a => 72, b => 291, p => true), (a => 73, b => 290, p => true), (a => 74, b => 289, p => true), (a => 75, b => 288, p => true), (a => 76, b => 287, p => true), (a => 77, b => 286, p => true), (a => 78, b => 285, p => true), (a => 79, b => 284, p => true), (a => 80, b => 283, p => true), (a => 81, b => 282, p => true), (a => 82, b => 281, p => true), (a => 83, b => 280, p => true), (a => 84, b => 279, p => true), (a => 85, b => 278, p => true), (a => 86, b => 277, p => true), (a => 87, b => 276, p => true), (a => 88, b => 275, p => true), (a => 89, b => 274, p => true), (a => 90, b => 273, p => true), (a => 91, b => 272, p => true), (a => 92, b => 271, p => true), (a => 93, b => 270, p => true), (a => 94, b => 269, p => true), (a => 95, b => 268, p => true), (a => 96, b => 267, p => true), (a => 97, b => 266, p => true), (a => 98, b => 265, p => true), (a => 99, b => 264, p => true), (a => 100, b => 263, p => true), (a => 101, b => 262, p => true), (a => 102, b => 261, p => true), (a => 103, b => 260, p => true), (a => 104, b => 259, p => true), (a => 105, b => 258, p => true), (a => 106, b => 257, p => true), (a => 107, b => 256, p => true), (a => 108, b => 255, p => true), (a => 109, b => 254, p => true), (a => 110, b => 253, p => true), (a => 111, b => 252, p => true), (a => 112, b => 251, p => true), (a => 113, b => 250, p => true), (a => 114, b => 249, p => true), (a => 115, b => 248, p => true), (a => 116, b => 247, p => true), (a => 117, b => 246, p => true), (a => 118, b => 245, p => true), (a => 119, b => 244, p => true), (a => 120, b => 243, p => true), (a => 121, b => 242, p => true), (a => 122, b => 241, p => true), (a => 123, b => 240, p => true), (a => 124, b => 239, p => true), (a => 125, b => 238, p => true), (a => 126, b => 237, p => true), (a => 127, b => 236, p => true), (a => 128, b => 235, p => true), (a => 129, b => 234, p => true), (a => 130, b => 233, p => true), (a => 131, b => 232, p => true), (a => 132, b => 231, p => true), (a => 133, b => 230, p => true), (a => 134, b => 229, p => true), (a => 135, b => 228, p => true), (a => 136, b => 227, p => true), (a => 137, b => 226, p => true), (a => 138, b => 225, p => true), (a => 139, b => 224, p => true), (a => 140, b => 223, p => true), (a => 141, b => 222, p => true), (a => 142, b => 221, p => true), (a => 143, b => 220, p => true), (a => 144, b => 219, p => true), (a => 145, b => 218, p => true), (a => 146, b => 217, p => true), (a => 147, b => 216, p => true), (a => 148, b => 215, p => true), (a => 149, b => 214, p => true), (a => 150, b => 213, p => true), (a => 151, b => 212, p => true), (a => 152, b => 211, p => true), (a => 153, b => 210, p => true), (a => 154, b => 209, p => true), (a => 155, b => 208, p => true), (a => 156, b => 207, p => true), (a => 157, b => 206, p => true), (a => 158, b => 205, p => true), (a => 159, b => 204, p => true), (a => 160, b => 203, p => true), (a => 161, b => 202, p => true), (a => 162, b => 201, p => true), (a => 163, b => 200, p => true), (a => 164, b => 199, p => true), (a => 165, b => 198, p => true), (a => 166, b => 197, p => true), (a => 167, b => 196, p => true), (a => 168, b => 195, p => true), (a => 169, b => 194, p => true), (a => 170, b => 193, p => true), (a => 171, b => 192, p => true), (a => 172, b => 191, p => true), (a => 173, b => 190, p => true), (a => 174, b => 189, p => true), (a => 175, b => 188, p => true), (a => 180, b => 187, p => true), (a => 181, b => 186, p => true), (a => 182, b => 185, p => true), (a => 183, b => 184, p => true)),
        ((a    => 2, b => 4, p => false), (a => 6, b => 8, p => false), (a => 10, b => 12, p => false), (a => 14, b => 176, p => false), (a => 3, b => 5, p => false), (a => 7, b => 9, p => false), (a => 11, b => 13, p => false), (a => 15, b => 177, p => false), (a => 0, b => 351, p => true), (a => 1, b => 350, p => true), (a => 16, b => 349, p => true), (a => 17, b => 348, p => true), (a => 18, b => 347, p => true), (a => 19, b => 346, p => true), (a => 20, b => 345, p => true), (a => 21, b => 344, p => true), (a => 22, b => 343, p => true), (a => 23, b => 342, p => true), (a => 24, b => 341, p => true), (a => 25, b => 340, p => true), (a => 26, b => 339, p => true), (a => 27, b => 338, p => true), (a => 28, b => 337, p => true), (a => 29, b => 336, p => true), (a => 30, b => 335, p => true), (a => 31, b => 334, p => true), (a => 32, b => 333, p => true), (a => 33, b => 332, p => true), (a => 34, b => 331, p => true), (a => 35, b => 330, p => true), (a => 36, b => 329, p => true), (a => 37, b => 328, p => true), (a => 38, b => 327, p => true), (a => 39, b => 326, p => true), (a => 40, b => 325, p => true), (a => 41, b => 324, p => true), (a => 42, b => 323, p => true), (a => 43, b => 322, p => true), (a => 44, b => 321, p => true), (a => 45, b => 320, p => true), (a => 46, b => 319, p => true), (a => 47, b => 318, p => true), (a => 48, b => 317, p => true), (a => 49, b => 316, p => true), (a => 50, b => 315, p => true), (a => 51, b => 314, p => true), (a => 52, b => 313, p => true), (a => 53, b => 312, p => true), (a => 54, b => 311, p => true), (a => 55, b => 310, p => true), (a => 56, b => 309, p => true), (a => 57, b => 308, p => true), (a => 58, b => 307, p => true), (a => 59, b => 306, p => true), (a => 60, b => 305, p => true), (a => 61, b => 304, p => true), (a => 62, b => 303, p => true), (a => 63, b => 302, p => true), (a => 64, b => 301, p => true), (a => 65, b => 300, p => true), (a => 66, b => 299, p => true), (a => 67, b => 298, p => true), (a => 68, b => 297, p => true), (a => 69, b => 296, p => true), (a => 70, b => 295, p => true), (a => 71, b => 294, p => true), (a => 72, b => 293, p => true), (a => 73, b => 292, p => true), (a => 74, b => 291, p => true), (a => 75, b => 290, p => true), (a => 76, b => 289, p => true), (a => 77, b => 288, p => true), (a => 78, b => 287, p => true), (a => 79, b => 286, p => true), (a => 80, b => 285, p => true), (a => 81, b => 284, p => true), (a => 82, b => 283, p => true), (a => 83, b => 282, p => true), (a => 84, b => 281, p => true), (a => 85, b => 280, p => true), (a => 86, b => 279, p => true), (a => 87, b => 278, p => true), (a => 88, b => 277, p => true), (a => 89, b => 276, p => true), (a => 90, b => 275, p => true), (a => 91, b => 274, p => true), (a => 92, b => 273, p => true), (a => 93, b => 272, p => true), (a => 94, b => 271, p => true), (a => 95, b => 270, p => true), (a => 96, b => 269, p => true), (a => 97, b => 268, p => true), (a => 98, b => 267, p => true), (a => 99, b => 266, p => true), (a => 100, b => 265, p => true), (a => 101, b => 264, p => true), (a => 102, b => 263, p => true), (a => 103, b => 262, p => true), (a => 104, b => 261, p => true), (a => 105, b => 260, p => true), (a => 106, b => 259, p => true), (a => 107, b => 258, p => true), (a => 108, b => 257, p => true), (a => 109, b => 256, p => true), (a => 110, b => 255, p => true), (a => 111, b => 254, p => true), (a => 112, b => 253, p => true), (a => 113, b => 252, p => true), (a => 114, b => 251, p => true), (a => 115, b => 250, p => true), (a => 116, b => 249, p => true), (a => 117, b => 248, p => true), (a => 118, b => 247, p => true), (a => 119, b => 246, p => true), (a => 120, b => 245, p => true), (a => 121, b => 244, p => true), (a => 122, b => 243, p => true), (a => 123, b => 242, p => true), (a => 124, b => 241, p => true), (a => 125, b => 240, p => true), (a => 126, b => 239, p => true), (a => 127, b => 238, p => true), (a => 128, b => 237, p => true), (a => 129, b => 236, p => true), (a => 130, b => 235, p => true), (a => 131, b => 234, p => true), (a => 132, b => 233, p => true), (a => 133, b => 232, p => true), (a => 134, b => 231, p => true), (a => 135, b => 230, p => true), (a => 136, b => 229, p => true), (a => 137, b => 228, p => true), (a => 138, b => 227, p => true), (a => 139, b => 226, p => true), (a => 140, b => 225, p => true), (a => 141, b => 224, p => true), (a => 142, b => 223, p => true), (a => 143, b => 222, p => true), (a => 144, b => 221, p => true), (a => 145, b => 220, p => true), (a => 146, b => 219, p => true), (a => 147, b => 218, p => true), (a => 148, b => 217, p => true), (a => 149, b => 216, p => true), (a => 150, b => 215, p => true), (a => 151, b => 214, p => true), (a => 152, b => 213, p => true), (a => 153, b => 212, p => true), (a => 154, b => 211, p => true), (a => 155, b => 210, p => true), (a => 156, b => 209, p => true), (a => 157, b => 208, p => true), (a => 158, b => 207, p => true), (a => 159, b => 206, p => true), (a => 160, b => 205, p => true), (a => 161, b => 204, p => true), (a => 162, b => 203, p => true), (a => 163, b => 202, p => true), (a => 164, b => 201, p => true), (a => 165, b => 200, p => true), (a => 166, b => 199, p => true), (a => 167, b => 198, p => true), (a => 168, b => 197, p => true), (a => 169, b => 196, p => true), (a => 170, b => 195, p => true), (a => 171, b => 194, p => true), (a => 172, b => 193, p => true), (a => 173, b => 192, p => true), (a => 174, b => 191, p => true), (a => 175, b => 190, p => true), (a => 178, b => 189, p => true), (a => 179, b => 188, p => true), (a => 180, b => 187, p => true), (a => 181, b => 186, p => true), (a => 182, b => 185, p => true), (a => 183, b => 184, p => true)),
        ((a    => 1, b => 2, p => false), (a => 3, b => 4, p => false), (a => 5, b => 6, p => false), (a => 7, b => 8, p => false), (a => 9, b => 10, p => false), (a => 11, b => 12, p => false), (a => 13, b => 14, p => false), (a => 15, b => 176, p => false), (a => 0, b => 351, p => true), (a => 16, b => 350, p => true), (a => 17, b => 349, p => true), (a => 18, b => 348, p => true), (a => 19, b => 347, p => true), (a => 20, b => 346, p => true), (a => 21, b => 345, p => true), (a => 22, b => 344, p => true), (a => 23, b => 343, p => true), (a => 24, b => 342, p => true), (a => 25, b => 341, p => true), (a => 26, b => 340, p => true), (a => 27, b => 339, p => true), (a => 28, b => 338, p => true), (a => 29, b => 337, p => true), (a => 30, b => 336, p => true), (a => 31, b => 335, p => true), (a => 32, b => 334, p => true), (a => 33, b => 333, p => true), (a => 34, b => 332, p => true), (a => 35, b => 331, p => true), (a => 36, b => 330, p => true), (a => 37, b => 329, p => true), (a => 38, b => 328, p => true), (a => 39, b => 327, p => true), (a => 40, b => 326, p => true), (a => 41, b => 325, p => true), (a => 42, b => 324, p => true), (a => 43, b => 323, p => true), (a => 44, b => 322, p => true), (a => 45, b => 321, p => true), (a => 46, b => 320, p => true), (a => 47, b => 319, p => true), (a => 48, b => 318, p => true), (a => 49, b => 317, p => true), (a => 50, b => 316, p => true), (a => 51, b => 315, p => true), (a => 52, b => 314, p => true), (a => 53, b => 313, p => true), (a => 54, b => 312, p => true), (a => 55, b => 311, p => true), (a => 56, b => 310, p => true), (a => 57, b => 309, p => true), (a => 58, b => 308, p => true), (a => 59, b => 307, p => true), (a => 60, b => 306, p => true), (a => 61, b => 305, p => true), (a => 62, b => 304, p => true), (a => 63, b => 303, p => true), (a => 64, b => 302, p => true), (a => 65, b => 301, p => true), (a => 66, b => 300, p => true), (a => 67, b => 299, p => true), (a => 68, b => 298, p => true), (a => 69, b => 297, p => true), (a => 70, b => 296, p => true), (a => 71, b => 295, p => true), (a => 72, b => 294, p => true), (a => 73, b => 293, p => true), (a => 74, b => 292, p => true), (a => 75, b => 291, p => true), (a => 76, b => 290, p => true), (a => 77, b => 289, p => true), (a => 78, b => 288, p => true), (a => 79, b => 287, p => true), (a => 80, b => 286, p => true), (a => 81, b => 285, p => true), (a => 82, b => 284, p => true), (a => 83, b => 283, p => true), (a => 84, b => 282, p => true), (a => 85, b => 281, p => true), (a => 86, b => 280, p => true), (a => 87, b => 279, p => true), (a => 88, b => 278, p => true), (a => 89, b => 277, p => true), (a => 90, b => 276, p => true), (a => 91, b => 275, p => true), (a => 92, b => 274, p => true), (a => 93, b => 273, p => true), (a => 94, b => 272, p => true), (a => 95, b => 271, p => true), (a => 96, b => 270, p => true), (a => 97, b => 269, p => true), (a => 98, b => 268, p => true), (a => 99, b => 267, p => true), (a => 100, b => 266, p => true), (a => 101, b => 265, p => true), (a => 102, b => 264, p => true), (a => 103, b => 263, p => true), (a => 104, b => 262, p => true), (a => 105, b => 261, p => true), (a => 106, b => 260, p => true), (a => 107, b => 259, p => true), (a => 108, b => 258, p => true), (a => 109, b => 257, p => true), (a => 110, b => 256, p => true), (a => 111, b => 255, p => true), (a => 112, b => 254, p => true), (a => 113, b => 253, p => true), (a => 114, b => 252, p => true), (a => 115, b => 251, p => true), (a => 116, b => 250, p => true), (a => 117, b => 249, p => true), (a => 118, b => 248, p => true), (a => 119, b => 247, p => true), (a => 120, b => 246, p => true), (a => 121, b => 245, p => true), (a => 122, b => 244, p => true), (a => 123, b => 243, p => true), (a => 124, b => 242, p => true), (a => 125, b => 241, p => true), (a => 126, b => 240, p => true), (a => 127, b => 239, p => true), (a => 128, b => 238, p => true), (a => 129, b => 237, p => true), (a => 130, b => 236, p => true), (a => 131, b => 235, p => true), (a => 132, b => 234, p => true), (a => 133, b => 233, p => true), (a => 134, b => 232, p => true), (a => 135, b => 231, p => true), (a => 136, b => 230, p => true), (a => 137, b => 229, p => true), (a => 138, b => 228, p => true), (a => 139, b => 227, p => true), (a => 140, b => 226, p => true), (a => 141, b => 225, p => true), (a => 142, b => 224, p => true), (a => 143, b => 223, p => true), (a => 144, b => 222, p => true), (a => 145, b => 221, p => true), (a => 146, b => 220, p => true), (a => 147, b => 219, p => true), (a => 148, b => 218, p => true), (a => 149, b => 217, p => true), (a => 150, b => 216, p => true), (a => 151, b => 215, p => true), (a => 152, b => 214, p => true), (a => 153, b => 213, p => true), (a => 154, b => 212, p => true), (a => 155, b => 211, p => true), (a => 156, b => 210, p => true), (a => 157, b => 209, p => true), (a => 158, b => 208, p => true), (a => 159, b => 207, p => true), (a => 160, b => 206, p => true), (a => 161, b => 205, p => true), (a => 162, b => 204, p => true), (a => 163, b => 203, p => true), (a => 164, b => 202, p => true), (a => 165, b => 201, p => true), (a => 166, b => 200, p => true), (a => 167, b => 199, p => true), (a => 168, b => 198, p => true), (a => 169, b => 197, p => true), (a => 170, b => 196, p => true), (a => 171, b => 195, p => true), (a => 172, b => 194, p => true), (a => 173, b => 193, p => true), (a => 174, b => 192, p => true), (a => 175, b => 191, p => true), (a => 177, b => 190, p => true), (a => 178, b => 189, p => true), (a => 179, b => 188, p => true), (a => 180, b => 187, p => true), (a => 181, b => 186, p => true), (a => 182, b => 185, p => true), (a => 183, b => 184, p => true))
        );


      when others => return empty_cfg;

    end case;
  end function get_cfg;

  function get_stg_off(depth : integer; D : integer; Off : integer) return stages_a is
    constant stage_a_d : stages_a := get_stg(352, D);
  begin
    return stage_a_d(Off to Off+depth-1);
  end function get_stg_off;

  function get_stg(I : integer; D : integer) return stages_a is
  begin
    case I is
      -- pipleline options for a total of 32 comparison stages
      -- 4 registers (D=4) is ok for implementing the whole sorting netwrok in the MSP FPGA
      when 352 =>
        case D is
          when 1 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, true);
                                        -- total number of registered stages: 1.
          when 2 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, true, false, false, false, false, false, false, false, false, false, false, false, false, false, false, false, true);
                                        -- total number of registered stages: 2.
          when 3 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, false, false, false, false, false, false, true, false, false, false, false, false, false, false, false, false, false, true, false, false, false, false, false, false, false, false, false, false, true);
                                        -- total number of registered stages: 3.
          when 4 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, false, false, false, false, true, false, false, false, false, false, false, false, true, false, false, false, false, false, false, false, true, false, false, false, false, false, false, false, true);
                                        -- total number of registered stages: 4.
          when 5 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, false, false, false, true, false, false, false, false, false, true, false, false, false, false, false, false, true, false, false, false, false, false, true, false, false, false, false, false, true);
                                        -- total number of registered stages: 5.
          when 6 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, false, false, true, false, false, false, false, true, false, false, false, false, false, true, false, false, false, false, true, false, false, false, false, true, false, false, false, false, true);
                                        -- total number of registered stages: 6.
          when 7 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, true, false, false, false, false, true, false, false, false, true, false, false, false, false, true, false, false, false, true, false, false, false, false, true, false, false, false, false, true);
                                        -- total number of registered stages: 7.
          when 8 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, true, false, false, false, true, false, false, false, true, false, false, false, true, false, false, false, true, false, false, false, true, false, false, false, true, false, false, false, true);
                                        -- total number of registered stages: 8.
          when 9 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, true, false, false, false, true, false, false, true, false, false, false, true, false, false, true, false, false, false, true, false, false, true, false, false, false, true, false, false, false, true);
                                        -- total number of registered stages: 9.
          when 10 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, false, true, false, false, true, false, false, true, false, false, true, false, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true);
                                        -- total number of registered stages: 10.
          when 11 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true, false, false, true);
                                        -- total number of registered stages: 11.
          when 12 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, false, false, true, false, false, true, false, true, false, false, true, false, false, true, false, true, false, false, true, false, false, true, false, true, false, false, true, false, false, true);
                                        -- total number of registered stages: 12.
          when 13 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, true, false, true, false, false, true, false, true, false, false, true, false, true, false, false, true, false, true, false, false, true, false, true, false, false, true, false, true, false, true);
                                        -- total number of registered stages: 13.
          when 14 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, true, false, true, false, true, false, false, true, false, true, false, true, false, false, true, false, true, false, true, false, true, false, false, true, false, true, false, true, false, true);
                                        -- total number of registered stages: 14.
          when 15 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true);
                                        -- total number of registered stages: 15.
          when 16 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true);
                                        -- total number of registered stages: 16.
          when 17 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true, false, true);
                                        -- total number of registered stages: 17.
          when 18 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (true, false, true, false, true, false, true, true, false, true, false, true, false, true, false, true, true, false, true, false, true, false, true, true, false, true, false, true, false, true, false, true);
                                        -- total number of registered stages: 18.
          when 19 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (true, false, true, false, true, true, false, true, false, true, true, false, true, false, true, true, false, true, false, true, true, false, true, false, true, true, false, true, false, true, false, true);
                                        -- total number of registered stages: 19.
          when 20 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (true, false, true, true, false, true, false, true, true, false, true, true, false, true, false, true, true, false, true, true, false, true, false, true, true, false, true, true, false, true, false, true);
                                        -- total number of registered stages: 20.
          when 21 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, false, true);
                                        -- total number of registered stages: 21.
          when 22 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, false, true, true, true, false, true, true, false, true, true, false, true, true, false, true, true, true);
                                        -- total number of registered stages: 22.
          when 23 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, false, true, true, true, false, true, true, false, true, true, true, false, true, true, false, true, true, true, false, true, true, false, true, true, true, false, true, true, true);
                                        -- total number of registered stages: 23.
          when 24 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, false, true, true, true, false, true, true, true, false, true, true, true, false, true, true, true, false, true, true, true, false, true, true, true, false, true, true, true, true);
                                        -- total number of registered stages: 24.
          when 25 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, false, true, true, true, true, false, true, true, true, false, true, true, true, true, false, true, true, true, false, true, true, true, true, false, true, true, true, true);
                                        -- total number of registered stages: 25.
          when 26 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, true, false, true, true, true, true, false, true, true, true, true, false, true, true, true, true, true, false, true, true, true, true, false, true, true, true, true, true);
                                        -- total number of registered stages: 26.
          when 27 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, true, true, false, true, true, true, true, true, false, true, true, true, true, true, true, false, true, true, true, true, true, false, true, true, true, true, true, true);
                                        -- total number of registered stages: 27.
          when 28 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, true, true, true, false, true, true, true, true, true, true, true, false, true, true, true, true, true, true, true, false, true, true, true, true, true, true, true, true);
                                        -- total number of registered stages: 28.
          when 29 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, true, true, true, true, true, true, false, true, true, true, true, true, true, true, true, true, true, false, true, true, true, true, true, true, true, true, true, true);
                                        -- total number of registered stages: 29.
          when 30 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, true, true, true, true, true, true, true, true, true, true, true, false, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true);
                                        -- total number of registered stages: 30.
          when 31 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (false, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true);
                                        -- total number of registered stages: 31.
          when 32 =>
                                        -- Registered stages configuration
                                        -- num -> |     0,     1,     2,     3,     4,     5,     6,     7,     8,     9,    10,    11,    12,    13,    14,    15,    16,    17,    18,    19,    20,    21,    22,    23,    24,    25,    26,    27,    28,    29,    30,    31|;
            return (true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true, true);
                                        -- total number of registered stages: 32.

          when others =>
            null;
        end case;

      when others => return (false, false);

    end case;
  end function get_stg;

  function to_array(data : std_logic_vector; N : integer) return muon_a is
    variable muon  : muon_a(0 to N - 1);
    variable left  : integer;
    variable right : integer;
  begin
    for i in muon'range loop
      left          := (i + 1) * in_word_w - 1;
      right         := i * in_word_w;
      muon(i).pt    := data(left - FLAGS_WIDTH - ROI_WIDTH downto right);
      muon(i).roi   := data(left - FLAGS_WIDTH downto right + PT_WIDTH);
      muon(i).flags := data(left downto right + PT_WIDTH + ROI_WIDTH);
    end loop;
    return muon;
  end to_array;

  function to_stdv(muon : muon_a; N : integer) return std_logic_vector is
    variable data  : std_logic_vector(N * out_word_w - 1 downto 0);
    variable left  : integer;
    variable right : integer;
  begin
    for i in muon'range loop
      left                                                          := (i + 1) * out_word_w - 1;
      right                                                         := i * out_word_w;
      data(left - IDX_WIDTH - FLAGS_WIDTH - ROI_WIDTH downto right) := muon(i).pt;
      data(left - IDX_WIDTH - FLAGS_WIDTH downto right + PT_WIDTH)  := muon(i).roi;
      data(left - IDX_WIDTH downto right + PT_WIDTH + ROI_WIDTH)    := muon(i).flags;
      data(left downto right + PT_WIDTH + ROI_WIDTH + FLAGS_WIDTH)  := muon(i).idx;
    end loop;
    return data;
  end to_stdv;

end package body csn_pkg;
