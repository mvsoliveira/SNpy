library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity compare_wrapper is

  port (
    ap_clk          : in  std_logic;
    ap_rst          : in  std_logic;
    ap_start        : in  std_logic;
    ap_done         : out std_logic;
    ap_idle         : out std_logic;
    ap_ready        : out std_logic;
    idata_0_pt_V    : in  std_logic_vector (3 downto 0);
    idata_1_pt_V    : in  std_logic_vector (3 downto 0);
    idata_2_pt_V    : in  std_logic_vector (3 downto 0);
    idata_3_pt_V    : in  std_logic_vector (3 downto 0);
    idata_4_pt_V    : in  std_logic_vector (3 downto 0);
    idata_5_pt_V    : in  std_logic_vector (3 downto 0);
    idata_6_pt_V    : in  std_logic_vector (3 downto 0);
    idata_7_pt_V    : in  std_logic_vector (3 downto 0);
    idata_8_pt_V    : in  std_logic_vector (3 downto 0);
    idata_9_pt_V    : in  std_logic_vector (3 downto 0);
    idata_10_pt_V   : in  std_logic_vector (3 downto 0);
    idata_11_pt_V   : in  std_logic_vector (3 downto 0);
    idata_12_pt_V   : in  std_logic_vector (3 downto 0);
    idata_13_pt_V   : in  std_logic_vector (3 downto 0);
    idata_14_pt_V   : in  std_logic_vector (3 downto 0);
    idata_15_pt_V   : in  std_logic_vector (3 downto 0);
    idata_16_pt_V   : in  std_logic_vector (3 downto 0);
    idata_17_pt_V   : in  std_logic_vector (3 downto 0);
    idata_18_pt_V   : in  std_logic_vector (3 downto 0);
    idata_19_pt_V   : in  std_logic_vector (3 downto 0);
    idata_20_pt_V   : in  std_logic_vector (3 downto 0);
    idata_21_pt_V   : in  std_logic_vector (3 downto 0);
    idata_22_pt_V   : in  std_logic_vector (3 downto 0);
    idata_23_pt_V   : in  std_logic_vector (3 downto 0);
    idata_24_pt_V   : in  std_logic_vector (3 downto 0);
    idata_25_pt_V   : in  std_logic_vector (3 downto 0);
    idata_26_pt_V   : in  std_logic_vector (3 downto 0);
    idata_27_pt_V   : in  std_logic_vector (3 downto 0);
    idata_28_pt_V   : in  std_logic_vector (3 downto 0);
    idata_29_pt_V   : in  std_logic_vector (3 downto 0);
    idata_30_pt_V   : in  std_logic_vector (3 downto 0);
    idata_31_pt_V   : in  std_logic_vector (3 downto 0);
    idata_32_pt_V   : in  std_logic_vector (3 downto 0);
    idata_33_pt_V   : in  std_logic_vector (3 downto 0);
    idata_34_pt_V   : in  std_logic_vector (3 downto 0);
    idata_35_pt_V   : in  std_logic_vector (3 downto 0);
    idata_36_pt_V   : in  std_logic_vector (3 downto 0);
    idata_37_pt_V   : in  std_logic_vector (3 downto 0);
    idata_38_pt_V   : in  std_logic_vector (3 downto 0);
    idata_39_pt_V   : in  std_logic_vector (3 downto 0);
    idata_40_pt_V   : in  std_logic_vector (3 downto 0);
    idata_41_pt_V   : in  std_logic_vector (3 downto 0);
    idata_42_pt_V   : in  std_logic_vector (3 downto 0);
    idata_43_pt_V   : in  std_logic_vector (3 downto 0);
    idata_44_pt_V   : in  std_logic_vector (3 downto 0);
    idata_45_pt_V   : in  std_logic_vector (3 downto 0);
    idata_46_pt_V   : in  std_logic_vector (3 downto 0);
    idata_47_pt_V   : in  std_logic_vector (3 downto 0);
    idata_48_pt_V   : in  std_logic_vector (3 downto 0);
    idata_49_pt_V   : in  std_logic_vector (3 downto 0);
    idata_50_pt_V   : in  std_logic_vector (3 downto 0);
    idata_51_pt_V   : in  std_logic_vector (3 downto 0);
    idata_52_pt_V   : in  std_logic_vector (3 downto 0);
    idata_53_pt_V   : in  std_logic_vector (3 downto 0);
    idata_54_pt_V   : in  std_logic_vector (3 downto 0);
    idata_55_pt_V   : in  std_logic_vector (3 downto 0);
    idata_56_pt_V   : in  std_logic_vector (3 downto 0);
    idata_57_pt_V   : in  std_logic_vector (3 downto 0);
    idata_58_pt_V   : in  std_logic_vector (3 downto 0);
    idata_59_pt_V   : in  std_logic_vector (3 downto 0);
    idata_60_pt_V   : in  std_logic_vector (3 downto 0);
    idata_61_pt_V   : in  std_logic_vector (3 downto 0);
    idata_62_pt_V   : in  std_logic_vector (3 downto 0);
    idata_63_pt_V   : in  std_logic_vector (3 downto 0);
    idata_64_pt_V   : in  std_logic_vector (3 downto 0);
    idata_65_pt_V   : in  std_logic_vector (3 downto 0);
    idata_66_pt_V   : in  std_logic_vector (3 downto 0);
    idata_67_pt_V   : in  std_logic_vector (3 downto 0);
    idata_68_pt_V   : in  std_logic_vector (3 downto 0);
    idata_69_pt_V   : in  std_logic_vector (3 downto 0);
    idata_70_pt_V   : in  std_logic_vector (3 downto 0);
    idata_71_pt_V   : in  std_logic_vector (3 downto 0);
    idata_72_pt_V   : in  std_logic_vector (3 downto 0);
    idata_73_pt_V   : in  std_logic_vector (3 downto 0);
    idata_74_pt_V   : in  std_logic_vector (3 downto 0);
    idata_75_pt_V   : in  std_logic_vector (3 downto 0);
    idata_76_pt_V   : in  std_logic_vector (3 downto 0);
    idata_77_pt_V   : in  std_logic_vector (3 downto 0);
    idata_78_pt_V   : in  std_logic_vector (3 downto 0);
    idata_79_pt_V   : in  std_logic_vector (3 downto 0);
    idata_80_pt_V   : in  std_logic_vector (3 downto 0);
    idata_81_pt_V   : in  std_logic_vector (3 downto 0);
    idata_82_pt_V   : in  std_logic_vector (3 downto 0);
    idata_83_pt_V   : in  std_logic_vector (3 downto 0);
    idata_84_pt_V   : in  std_logic_vector (3 downto 0);
    idata_85_pt_V   : in  std_logic_vector (3 downto 0);
    idata_86_pt_V   : in  std_logic_vector (3 downto 0);
    idata_87_pt_V   : in  std_logic_vector (3 downto 0);
    idata_88_pt_V   : in  std_logic_vector (3 downto 0);
    idata_89_pt_V   : in  std_logic_vector (3 downto 0);
    idata_90_pt_V   : in  std_logic_vector (3 downto 0);
    idata_91_pt_V   : in  std_logic_vector (3 downto 0);
    idata_92_pt_V   : in  std_logic_vector (3 downto 0);
    idata_93_pt_V   : in  std_logic_vector (3 downto 0);
    idata_94_pt_V   : in  std_logic_vector (3 downto 0);
    idata_95_pt_V   : in  std_logic_vector (3 downto 0);
    idata_96_pt_V   : in  std_logic_vector (3 downto 0);
    idata_97_pt_V   : in  std_logic_vector (3 downto 0);
    idata_98_pt_V   : in  std_logic_vector (3 downto 0);
    idata_99_pt_V   : in  std_logic_vector (3 downto 0);
    idata_100_pt_V  : in  std_logic_vector (3 downto 0);
    idata_101_pt_V  : in  std_logic_vector (3 downto 0);
    idata_102_pt_V  : in  std_logic_vector (3 downto 0);
    idata_103_pt_V  : in  std_logic_vector (3 downto 0);
    idata_104_pt_V  : in  std_logic_vector (3 downto 0);
    idata_105_pt_V  : in  std_logic_vector (3 downto 0);
    idata_106_pt_V  : in  std_logic_vector (3 downto 0);
    idata_107_pt_V  : in  std_logic_vector (3 downto 0);
    idata_108_pt_V  : in  std_logic_vector (3 downto 0);
    idata_109_pt_V  : in  std_logic_vector (3 downto 0);
    idata_110_pt_V  : in  std_logic_vector (3 downto 0);
    idata_111_pt_V  : in  std_logic_vector (3 downto 0);
    idata_112_pt_V  : in  std_logic_vector (3 downto 0);
    idata_113_pt_V  : in  std_logic_vector (3 downto 0);
    idata_114_pt_V  : in  std_logic_vector (3 downto 0);
    idata_115_pt_V  : in  std_logic_vector (3 downto 0);
    idata_116_pt_V  : in  std_logic_vector (3 downto 0);
    idata_117_pt_V  : in  std_logic_vector (3 downto 0);
    idata_118_pt_V  : in  std_logic_vector (3 downto 0);
    idata_119_pt_V  : in  std_logic_vector (3 downto 0);
    idata_120_pt_V  : in  std_logic_vector (3 downto 0);
    idata_121_pt_V  : in  std_logic_vector (3 downto 0);
    idata_122_pt_V  : in  std_logic_vector (3 downto 0);
    idata_123_pt_V  : in  std_logic_vector (3 downto 0);
    idata_124_pt_V  : in  std_logic_vector (3 downto 0);
    idata_125_pt_V  : in  std_logic_vector (3 downto 0);
    idata_126_pt_V  : in  std_logic_vector (3 downto 0);
    idata_127_pt_V  : in  std_logic_vector (3 downto 0);
    idata_128_pt_V  : in  std_logic_vector (3 downto 0);
    idata_129_pt_V  : in  std_logic_vector (3 downto 0);
    idata_130_pt_V  : in  std_logic_vector (3 downto 0);
    idata_131_pt_V  : in  std_logic_vector (3 downto 0);
    idata_132_pt_V  : in  std_logic_vector (3 downto 0);
    idata_133_pt_V  : in  std_logic_vector (3 downto 0);
    idata_134_pt_V  : in  std_logic_vector (3 downto 0);
    idata_135_pt_V  : in  std_logic_vector (3 downto 0);
    idata_136_pt_V  : in  std_logic_vector (3 downto 0);
    idata_137_pt_V  : in  std_logic_vector (3 downto 0);
    idata_138_pt_V  : in  std_logic_vector (3 downto 0);
    idata_139_pt_V  : in  std_logic_vector (3 downto 0);
    idata_140_pt_V  : in  std_logic_vector (3 downto 0);
    idata_141_pt_V  : in  std_logic_vector (3 downto 0);
    idata_142_pt_V  : in  std_logic_vector (3 downto 0);
    idata_143_pt_V  : in  std_logic_vector (3 downto 0);
    idata_144_pt_V  : in  std_logic_vector (3 downto 0);
    idata_145_pt_V  : in  std_logic_vector (3 downto 0);
    idata_146_pt_V  : in  std_logic_vector (3 downto 0);
    idata_147_pt_V  : in  std_logic_vector (3 downto 0);
    idata_148_pt_V  : in  std_logic_vector (3 downto 0);
    idata_149_pt_V  : in  std_logic_vector (3 downto 0);
    idata_150_pt_V  : in  std_logic_vector (3 downto 0);
    idata_151_pt_V  : in  std_logic_vector (3 downto 0);
    idata_152_pt_V  : in  std_logic_vector (3 downto 0);
    idata_153_pt_V  : in  std_logic_vector (3 downto 0);
    idata_154_pt_V  : in  std_logic_vector (3 downto 0);
    idata_155_pt_V  : in  std_logic_vector (3 downto 0);
    idata_156_pt_V  : in  std_logic_vector (3 downto 0);
    idata_157_pt_V  : in  std_logic_vector (3 downto 0);
    idata_158_pt_V  : in  std_logic_vector (3 downto 0);
    idata_159_pt_V  : in  std_logic_vector (3 downto 0);
    idata_160_pt_V  : in  std_logic_vector (3 downto 0);
    idata_161_pt_V  : in  std_logic_vector (3 downto 0);
    idata_162_pt_V  : in  std_logic_vector (3 downto 0);
    idata_163_pt_V  : in  std_logic_vector (3 downto 0);
    idata_164_pt_V  : in  std_logic_vector (3 downto 0);
    idata_165_pt_V  : in  std_logic_vector (3 downto 0);
    idata_166_pt_V  : in  std_logic_vector (3 downto 0);
    idata_167_pt_V  : in  std_logic_vector (3 downto 0);
    idata_168_pt_V  : in  std_logic_vector (3 downto 0);
    idata_169_pt_V  : in  std_logic_vector (3 downto 0);
    idata_170_pt_V  : in  std_logic_vector (3 downto 0);
    idata_171_pt_V  : in  std_logic_vector (3 downto 0);
    idata_172_pt_V  : in  std_logic_vector (3 downto 0);
    idata_173_pt_V  : in  std_logic_vector (3 downto 0);
    idata_174_pt_V  : in  std_logic_vector (3 downto 0);
    idata_175_pt_V  : in  std_logic_vector (3 downto 0);
    idata_176_pt_V  : in  std_logic_vector (3 downto 0);
    idata_177_pt_V  : in  std_logic_vector (3 downto 0);
    idata_178_pt_V  : in  std_logic_vector (3 downto 0);
    idata_179_pt_V  : in  std_logic_vector (3 downto 0);
    idata_180_pt_V  : in  std_logic_vector (3 downto 0);
    idata_181_pt_V  : in  std_logic_vector (3 downto 0);
    idata_182_pt_V  : in  std_logic_vector (3 downto 0);
    idata_183_pt_V  : in  std_logic_vector (3 downto 0);
    idata_184_pt_V  : in  std_logic_vector (3 downto 0);
    idata_185_pt_V  : in  std_logic_vector (3 downto 0);
    idata_186_pt_V  : in  std_logic_vector (3 downto 0);
    idata_187_pt_V  : in  std_logic_vector (3 downto 0);
    idata_188_pt_V  : in  std_logic_vector (3 downto 0);
    idata_189_pt_V  : in  std_logic_vector (3 downto 0);
    idata_190_pt_V  : in  std_logic_vector (3 downto 0);
    idata_191_pt_V  : in  std_logic_vector (3 downto 0);
    idata_192_pt_V  : in  std_logic_vector (3 downto 0);
    idata_193_pt_V  : in  std_logic_vector (3 downto 0);
    idata_194_pt_V  : in  std_logic_vector (3 downto 0);
    idata_195_pt_V  : in  std_logic_vector (3 downto 0);
    idata_196_pt_V  : in  std_logic_vector (3 downto 0);
    idata_197_pt_V  : in  std_logic_vector (3 downto 0);
    idata_198_pt_V  : in  std_logic_vector (3 downto 0);
    idata_199_pt_V  : in  std_logic_vector (3 downto 0);
    idata_200_pt_V  : in  std_logic_vector (3 downto 0);
    idata_201_pt_V  : in  std_logic_vector (3 downto 0);
    idata_202_pt_V  : in  std_logic_vector (3 downto 0);
    idata_203_pt_V  : in  std_logic_vector (3 downto 0);
    idata_204_pt_V  : in  std_logic_vector (3 downto 0);
    idata_205_pt_V  : in  std_logic_vector (3 downto 0);
    idata_206_pt_V  : in  std_logic_vector (3 downto 0);
    idata_207_pt_V  : in  std_logic_vector (3 downto 0);
    idata_208_pt_V  : in  std_logic_vector (3 downto 0);
    idata_209_pt_V  : in  std_logic_vector (3 downto 0);
    idata_210_pt_V  : in  std_logic_vector (3 downto 0);
    idata_211_pt_V  : in  std_logic_vector (3 downto 0);
    idata_212_pt_V  : in  std_logic_vector (3 downto 0);
    idata_213_pt_V  : in  std_logic_vector (3 downto 0);
    idata_214_pt_V  : in  std_logic_vector (3 downto 0);
    idata_215_pt_V  : in  std_logic_vector (3 downto 0);
    idata_216_pt_V  : in  std_logic_vector (3 downto 0);
    idata_217_pt_V  : in  std_logic_vector (3 downto 0);
    idata_218_pt_V  : in  std_logic_vector (3 downto 0);
    idata_219_pt_V  : in  std_logic_vector (3 downto 0);
    idata_220_pt_V  : in  std_logic_vector (3 downto 0);
    idata_221_pt_V  : in  std_logic_vector (3 downto 0);
    idata_222_pt_V  : in  std_logic_vector (3 downto 0);
    idata_223_pt_V  : in  std_logic_vector (3 downto 0);
    idata_224_pt_V  : in  std_logic_vector (3 downto 0);
    idata_225_pt_V  : in  std_logic_vector (3 downto 0);
    idata_226_pt_V  : in  std_logic_vector (3 downto 0);
    idata_227_pt_V  : in  std_logic_vector (3 downto 0);
    idata_228_pt_V  : in  std_logic_vector (3 downto 0);
    idata_229_pt_V  : in  std_logic_vector (3 downto 0);
    idata_230_pt_V  : in  std_logic_vector (3 downto 0);
    idata_231_pt_V  : in  std_logic_vector (3 downto 0);
    idata_232_pt_V  : in  std_logic_vector (3 downto 0);
    idata_233_pt_V  : in  std_logic_vector (3 downto 0);
    idata_234_pt_V  : in  std_logic_vector (3 downto 0);
    idata_235_pt_V  : in  std_logic_vector (3 downto 0);
    idata_236_pt_V  : in  std_logic_vector (3 downto 0);
    idata_237_pt_V  : in  std_logic_vector (3 downto 0);
    idata_238_pt_V  : in  std_logic_vector (3 downto 0);
    idata_239_pt_V  : in  std_logic_vector (3 downto 0);
    idata_240_pt_V  : in  std_logic_vector (3 downto 0);
    idata_241_pt_V  : in  std_logic_vector (3 downto 0);
    idata_242_pt_V  : in  std_logic_vector (3 downto 0);
    idata_243_pt_V  : in  std_logic_vector (3 downto 0);
    idata_244_pt_V  : in  std_logic_vector (3 downto 0);
    idata_245_pt_V  : in  std_logic_vector (3 downto 0);
    idata_246_pt_V  : in  std_logic_vector (3 downto 0);
    idata_247_pt_V  : in  std_logic_vector (3 downto 0);
    idata_248_pt_V  : in  std_logic_vector (3 downto 0);
    idata_249_pt_V  : in  std_logic_vector (3 downto 0);
    idata_250_pt_V  : in  std_logic_vector (3 downto 0);
    idata_251_pt_V  : in  std_logic_vector (3 downto 0);
    idata_252_pt_V  : in  std_logic_vector (3 downto 0);
    idata_253_pt_V  : in  std_logic_vector (3 downto 0);
    idata_254_pt_V  : in  std_logic_vector (3 downto 0);
    idata_255_pt_V  : in  std_logic_vector (3 downto 0);
    idata_256_pt_V  : in  std_logic_vector (3 downto 0);
    idata_257_pt_V  : in  std_logic_vector (3 downto 0);
    idata_258_pt_V  : in  std_logic_vector (3 downto 0);
    idata_259_pt_V  : in  std_logic_vector (3 downto 0);
    idata_260_pt_V  : in  std_logic_vector (3 downto 0);
    idata_261_pt_V  : in  std_logic_vector (3 downto 0);
    idata_262_pt_V  : in  std_logic_vector (3 downto 0);
    idata_263_pt_V  : in  std_logic_vector (3 downto 0);
    idata_264_pt_V  : in  std_logic_vector (3 downto 0);
    idata_265_pt_V  : in  std_logic_vector (3 downto 0);
    idata_266_pt_V  : in  std_logic_vector (3 downto 0);
    idata_267_pt_V  : in  std_logic_vector (3 downto 0);
    idata_268_pt_V  : in  std_logic_vector (3 downto 0);
    idata_269_pt_V  : in  std_logic_vector (3 downto 0);
    idata_270_pt_V  : in  std_logic_vector (3 downto 0);
    idata_271_pt_V  : in  std_logic_vector (3 downto 0);
    idata_272_pt_V  : in  std_logic_vector (3 downto 0);
    idata_273_pt_V  : in  std_logic_vector (3 downto 0);
    idata_274_pt_V  : in  std_logic_vector (3 downto 0);
    idata_275_pt_V  : in  std_logic_vector (3 downto 0);
    idata_276_pt_V  : in  std_logic_vector (3 downto 0);
    idata_277_pt_V  : in  std_logic_vector (3 downto 0);
    idata_278_pt_V  : in  std_logic_vector (3 downto 0);
    idata_279_pt_V  : in  std_logic_vector (3 downto 0);
    idata_280_pt_V  : in  std_logic_vector (3 downto 0);
    idata_281_pt_V  : in  std_logic_vector (3 downto 0);
    idata_282_pt_V  : in  std_logic_vector (3 downto 0);
    idata_283_pt_V  : in  std_logic_vector (3 downto 0);
    idata_284_pt_V  : in  std_logic_vector (3 downto 0);
    idata_285_pt_V  : in  std_logic_vector (3 downto 0);
    idata_286_pt_V  : in  std_logic_vector (3 downto 0);
    idata_287_pt_V  : in  std_logic_vector (3 downto 0);
    idata_288_pt_V  : in  std_logic_vector (3 downto 0);
    idata_289_pt_V  : in  std_logic_vector (3 downto 0);
    idata_290_pt_V  : in  std_logic_vector (3 downto 0);
    idata_291_pt_V  : in  std_logic_vector (3 downto 0);
    idata_292_pt_V  : in  std_logic_vector (3 downto 0);
    idata_293_pt_V  : in  std_logic_vector (3 downto 0);
    idata_294_pt_V  : in  std_logic_vector (3 downto 0);
    idata_295_pt_V  : in  std_logic_vector (3 downto 0);
    idata_296_pt_V  : in  std_logic_vector (3 downto 0);
    idata_297_pt_V  : in  std_logic_vector (3 downto 0);
    idata_298_pt_V  : in  std_logic_vector (3 downto 0);
    idata_299_pt_V  : in  std_logic_vector (3 downto 0);
    idata_300_pt_V  : in  std_logic_vector (3 downto 0);
    idata_301_pt_V  : in  std_logic_vector (3 downto 0);
    idata_302_pt_V  : in  std_logic_vector (3 downto 0);
    idata_303_pt_V  : in  std_logic_vector (3 downto 0);
    idata_304_pt_V  : in  std_logic_vector (3 downto 0);
    idata_305_pt_V  : in  std_logic_vector (3 downto 0);
    idata_306_pt_V  : in  std_logic_vector (3 downto 0);
    idata_307_pt_V  : in  std_logic_vector (3 downto 0);
    idata_308_pt_V  : in  std_logic_vector (3 downto 0);
    idata_309_pt_V  : in  std_logic_vector (3 downto 0);
    idata_310_pt_V  : in  std_logic_vector (3 downto 0);
    idata_311_pt_V  : in  std_logic_vector (3 downto 0);
    idata_312_pt_V  : in  std_logic_vector (3 downto 0);
    idata_313_pt_V  : in  std_logic_vector (3 downto 0);
    idata_314_pt_V  : in  std_logic_vector (3 downto 0);
    idata_315_pt_V  : in  std_logic_vector (3 downto 0);
    idata_316_pt_V  : in  std_logic_vector (3 downto 0);
    idata_317_pt_V  : in  std_logic_vector (3 downto 0);
    idata_318_pt_V  : in  std_logic_vector (3 downto 0);
    idata_319_pt_V  : in  std_logic_vector (3 downto 0);
    idata_320_pt_V  : in  std_logic_vector (3 downto 0);
    idata_321_pt_V  : in  std_logic_vector (3 downto 0);
    idata_322_pt_V  : in  std_logic_vector (3 downto 0);
    idata_323_pt_V  : in  std_logic_vector (3 downto 0);
    idata_324_pt_V  : in  std_logic_vector (3 downto 0);
    idata_325_pt_V  : in  std_logic_vector (3 downto 0);
    idata_326_pt_V  : in  std_logic_vector (3 downto 0);
    idata_327_pt_V  : in  std_logic_vector (3 downto 0);
    idata_328_pt_V  : in  std_logic_vector (3 downto 0);
    idata_329_pt_V  : in  std_logic_vector (3 downto 0);
    idata_330_pt_V  : in  std_logic_vector (3 downto 0);
    idata_331_pt_V  : in  std_logic_vector (3 downto 0);
    idata_332_pt_V  : in  std_logic_vector (3 downto 0);
    idata_333_pt_V  : in  std_logic_vector (3 downto 0);
    idata_334_pt_V  : in  std_logic_vector (3 downto 0);
    idata_335_pt_V  : in  std_logic_vector (3 downto 0);
    idata_336_pt_V  : in  std_logic_vector (3 downto 0);
    idata_337_pt_V  : in  std_logic_vector (3 downto 0);
    idata_338_pt_V  : in  std_logic_vector (3 downto 0);
    idata_339_pt_V  : in  std_logic_vector (3 downto 0);
    idata_340_pt_V  : in  std_logic_vector (3 downto 0);
    idata_341_pt_V  : in  std_logic_vector (3 downto 0);
    idata_342_pt_V  : in  std_logic_vector (3 downto 0);
    idata_343_pt_V  : in  std_logic_vector (3 downto 0);
    idata_344_pt_V  : in  std_logic_vector (3 downto 0);
    idata_345_pt_V  : in  std_logic_vector (3 downto 0);
    idata_346_pt_V  : in  std_logic_vector (3 downto 0);
    idata_347_pt_V  : in  std_logic_vector (3 downto 0);
    idata_348_pt_V  : in  std_logic_vector (3 downto 0);
    idata_349_pt_V  : in  std_logic_vector (3 downto 0);
    idata_350_pt_V  : in  std_logic_vector (3 downto 0);
    idata_351_pt_V  : in  std_logic_vector (3 downto 0);
    idata_0_roi_V   : in  std_logic_vector (7 downto 0);
    idata_1_roi_V   : in  std_logic_vector (7 downto 0);
    idata_2_roi_V   : in  std_logic_vector (7 downto 0);
    idata_3_roi_V   : in  std_logic_vector (7 downto 0);
    idata_4_roi_V   : in  std_logic_vector (7 downto 0);
    idata_5_roi_V   : in  std_logic_vector (7 downto 0);
    idata_6_roi_V   : in  std_logic_vector (7 downto 0);
    idata_7_roi_V   : in  std_logic_vector (7 downto 0);
    idata_8_roi_V   : in  std_logic_vector (7 downto 0);
    idata_9_roi_V   : in  std_logic_vector (7 downto 0);
    idata_10_roi_V  : in  std_logic_vector (7 downto 0);
    idata_11_roi_V  : in  std_logic_vector (7 downto 0);
    idata_12_roi_V  : in  std_logic_vector (7 downto 0);
    idata_13_roi_V  : in  std_logic_vector (7 downto 0);
    idata_14_roi_V  : in  std_logic_vector (7 downto 0);
    idata_15_roi_V  : in  std_logic_vector (7 downto 0);
    idata_16_roi_V  : in  std_logic_vector (7 downto 0);
    idata_17_roi_V  : in  std_logic_vector (7 downto 0);
    idata_18_roi_V  : in  std_logic_vector (7 downto 0);
    idata_19_roi_V  : in  std_logic_vector (7 downto 0);
    idata_20_roi_V  : in  std_logic_vector (7 downto 0);
    idata_21_roi_V  : in  std_logic_vector (7 downto 0);
    idata_22_roi_V  : in  std_logic_vector (7 downto 0);
    idata_23_roi_V  : in  std_logic_vector (7 downto 0);
    idata_24_roi_V  : in  std_logic_vector (7 downto 0);
    idata_25_roi_V  : in  std_logic_vector (7 downto 0);
    idata_26_roi_V  : in  std_logic_vector (7 downto 0);
    idata_27_roi_V  : in  std_logic_vector (7 downto 0);
    idata_28_roi_V  : in  std_logic_vector (7 downto 0);
    idata_29_roi_V  : in  std_logic_vector (7 downto 0);
    idata_30_roi_V  : in  std_logic_vector (7 downto 0);
    idata_31_roi_V  : in  std_logic_vector (7 downto 0);
    idata_32_roi_V  : in  std_logic_vector (7 downto 0);
    idata_33_roi_V  : in  std_logic_vector (7 downto 0);
    idata_34_roi_V  : in  std_logic_vector (7 downto 0);
    idata_35_roi_V  : in  std_logic_vector (7 downto 0);
    idata_36_roi_V  : in  std_logic_vector (7 downto 0);
    idata_37_roi_V  : in  std_logic_vector (7 downto 0);
    idata_38_roi_V  : in  std_logic_vector (7 downto 0);
    idata_39_roi_V  : in  std_logic_vector (7 downto 0);
    idata_40_roi_V  : in  std_logic_vector (7 downto 0);
    idata_41_roi_V  : in  std_logic_vector (7 downto 0);
    idata_42_roi_V  : in  std_logic_vector (7 downto 0);
    idata_43_roi_V  : in  std_logic_vector (7 downto 0);
    idata_44_roi_V  : in  std_logic_vector (7 downto 0);
    idata_45_roi_V  : in  std_logic_vector (7 downto 0);
    idata_46_roi_V  : in  std_logic_vector (7 downto 0);
    idata_47_roi_V  : in  std_logic_vector (7 downto 0);
    idata_48_roi_V  : in  std_logic_vector (7 downto 0);
    idata_49_roi_V  : in  std_logic_vector (7 downto 0);
    idata_50_roi_V  : in  std_logic_vector (7 downto 0);
    idata_51_roi_V  : in  std_logic_vector (7 downto 0);
    idata_52_roi_V  : in  std_logic_vector (7 downto 0);
    idata_53_roi_V  : in  std_logic_vector (7 downto 0);
    idata_54_roi_V  : in  std_logic_vector (7 downto 0);
    idata_55_roi_V  : in  std_logic_vector (7 downto 0);
    idata_56_roi_V  : in  std_logic_vector (7 downto 0);
    idata_57_roi_V  : in  std_logic_vector (7 downto 0);
    idata_58_roi_V  : in  std_logic_vector (7 downto 0);
    idata_59_roi_V  : in  std_logic_vector (7 downto 0);
    idata_60_roi_V  : in  std_logic_vector (7 downto 0);
    idata_61_roi_V  : in  std_logic_vector (7 downto 0);
    idata_62_roi_V  : in  std_logic_vector (7 downto 0);
    idata_63_roi_V  : in  std_logic_vector (7 downto 0);
    idata_64_roi_V  : in  std_logic_vector (7 downto 0);
    idata_65_roi_V  : in  std_logic_vector (7 downto 0);
    idata_66_roi_V  : in  std_logic_vector (7 downto 0);
    idata_67_roi_V  : in  std_logic_vector (7 downto 0);
    idata_68_roi_V  : in  std_logic_vector (7 downto 0);
    idata_69_roi_V  : in  std_logic_vector (7 downto 0);
    idata_70_roi_V  : in  std_logic_vector (7 downto 0);
    idata_71_roi_V  : in  std_logic_vector (7 downto 0);
    idata_72_roi_V  : in  std_logic_vector (7 downto 0);
    idata_73_roi_V  : in  std_logic_vector (7 downto 0);
    idata_74_roi_V  : in  std_logic_vector (7 downto 0);
    idata_75_roi_V  : in  std_logic_vector (7 downto 0);
    idata_76_roi_V  : in  std_logic_vector (7 downto 0);
    idata_77_roi_V  : in  std_logic_vector (7 downto 0);
    idata_78_roi_V  : in  std_logic_vector (7 downto 0);
    idata_79_roi_V  : in  std_logic_vector (7 downto 0);
    idata_80_roi_V  : in  std_logic_vector (7 downto 0);
    idata_81_roi_V  : in  std_logic_vector (7 downto 0);
    idata_82_roi_V  : in  std_logic_vector (7 downto 0);
    idata_83_roi_V  : in  std_logic_vector (7 downto 0);
    idata_84_roi_V  : in  std_logic_vector (7 downto 0);
    idata_85_roi_V  : in  std_logic_vector (7 downto 0);
    idata_86_roi_V  : in  std_logic_vector (7 downto 0);
    idata_87_roi_V  : in  std_logic_vector (7 downto 0);
    idata_88_roi_V  : in  std_logic_vector (7 downto 0);
    idata_89_roi_V  : in  std_logic_vector (7 downto 0);
    idata_90_roi_V  : in  std_logic_vector (7 downto 0);
    idata_91_roi_V  : in  std_logic_vector (7 downto 0);
    idata_92_roi_V  : in  std_logic_vector (7 downto 0);
    idata_93_roi_V  : in  std_logic_vector (7 downto 0);
    idata_94_roi_V  : in  std_logic_vector (7 downto 0);
    idata_95_roi_V  : in  std_logic_vector (7 downto 0);
    idata_96_roi_V  : in  std_logic_vector (7 downto 0);
    idata_97_roi_V  : in  std_logic_vector (7 downto 0);
    idata_98_roi_V  : in  std_logic_vector (7 downto 0);
    idata_99_roi_V  : in  std_logic_vector (7 downto 0);
    idata_100_roi_V : in  std_logic_vector (7 downto 0);
    idata_101_roi_V : in  std_logic_vector (7 downto 0);
    idata_102_roi_V : in  std_logic_vector (7 downto 0);
    idata_103_roi_V : in  std_logic_vector (7 downto 0);
    idata_104_roi_V : in  std_logic_vector (7 downto 0);
    idata_105_roi_V : in  std_logic_vector (7 downto 0);
    idata_106_roi_V : in  std_logic_vector (7 downto 0);
    idata_107_roi_V : in  std_logic_vector (7 downto 0);
    idata_108_roi_V : in  std_logic_vector (7 downto 0);
    idata_109_roi_V : in  std_logic_vector (7 downto 0);
    idata_110_roi_V : in  std_logic_vector (7 downto 0);
    idata_111_roi_V : in  std_logic_vector (7 downto 0);
    idata_112_roi_V : in  std_logic_vector (7 downto 0);
    idata_113_roi_V : in  std_logic_vector (7 downto 0);
    idata_114_roi_V : in  std_logic_vector (7 downto 0);
    idata_115_roi_V : in  std_logic_vector (7 downto 0);
    idata_116_roi_V : in  std_logic_vector (7 downto 0);
    idata_117_roi_V : in  std_logic_vector (7 downto 0);
    idata_118_roi_V : in  std_logic_vector (7 downto 0);
    idata_119_roi_V : in  std_logic_vector (7 downto 0);
    idata_120_roi_V : in  std_logic_vector (7 downto 0);
    idata_121_roi_V : in  std_logic_vector (7 downto 0);
    idata_122_roi_V : in  std_logic_vector (7 downto 0);
    idata_123_roi_V : in  std_logic_vector (7 downto 0);
    idata_124_roi_V : in  std_logic_vector (7 downto 0);
    idata_125_roi_V : in  std_logic_vector (7 downto 0);
    idata_126_roi_V : in  std_logic_vector (7 downto 0);
    idata_127_roi_V : in  std_logic_vector (7 downto 0);
    idata_128_roi_V : in  std_logic_vector (7 downto 0);
    idata_129_roi_V : in  std_logic_vector (7 downto 0);
    idata_130_roi_V : in  std_logic_vector (7 downto 0);
    idata_131_roi_V : in  std_logic_vector (7 downto 0);
    idata_132_roi_V : in  std_logic_vector (7 downto 0);
    idata_133_roi_V : in  std_logic_vector (7 downto 0);
    idata_134_roi_V : in  std_logic_vector (7 downto 0);
    idata_135_roi_V : in  std_logic_vector (7 downto 0);
    idata_136_roi_V : in  std_logic_vector (7 downto 0);
    idata_137_roi_V : in  std_logic_vector (7 downto 0);
    idata_138_roi_V : in  std_logic_vector (7 downto 0);
    idata_139_roi_V : in  std_logic_vector (7 downto 0);
    idata_140_roi_V : in  std_logic_vector (7 downto 0);
    idata_141_roi_V : in  std_logic_vector (7 downto 0);
    idata_142_roi_V : in  std_logic_vector (7 downto 0);
    idata_143_roi_V : in  std_logic_vector (7 downto 0);
    idata_144_roi_V : in  std_logic_vector (7 downto 0);
    idata_145_roi_V : in  std_logic_vector (7 downto 0);
    idata_146_roi_V : in  std_logic_vector (7 downto 0);
    idata_147_roi_V : in  std_logic_vector (7 downto 0);
    idata_148_roi_V : in  std_logic_vector (7 downto 0);
    idata_149_roi_V : in  std_logic_vector (7 downto 0);
    idata_150_roi_V : in  std_logic_vector (7 downto 0);
    idata_151_roi_V : in  std_logic_vector (7 downto 0);
    idata_152_roi_V : in  std_logic_vector (7 downto 0);
    idata_153_roi_V : in  std_logic_vector (7 downto 0);
    idata_154_roi_V : in  std_logic_vector (7 downto 0);
    idata_155_roi_V : in  std_logic_vector (7 downto 0);
    idata_156_roi_V : in  std_logic_vector (7 downto 0);
    idata_157_roi_V : in  std_logic_vector (7 downto 0);
    idata_158_roi_V : in  std_logic_vector (7 downto 0);
    idata_159_roi_V : in  std_logic_vector (7 downto 0);
    idata_160_roi_V : in  std_logic_vector (7 downto 0);
    idata_161_roi_V : in  std_logic_vector (7 downto 0);
    idata_162_roi_V : in  std_logic_vector (7 downto 0);
    idata_163_roi_V : in  std_logic_vector (7 downto 0);
    idata_164_roi_V : in  std_logic_vector (7 downto 0);
    idata_165_roi_V : in  std_logic_vector (7 downto 0);
    idata_166_roi_V : in  std_logic_vector (7 downto 0);
    idata_167_roi_V : in  std_logic_vector (7 downto 0);
    idata_168_roi_V : in  std_logic_vector (7 downto 0);
    idata_169_roi_V : in  std_logic_vector (7 downto 0);
    idata_170_roi_V : in  std_logic_vector (7 downto 0);
    idata_171_roi_V : in  std_logic_vector (7 downto 0);
    idata_172_roi_V : in  std_logic_vector (7 downto 0);
    idata_173_roi_V : in  std_logic_vector (7 downto 0);
    idata_174_roi_V : in  std_logic_vector (7 downto 0);
    idata_175_roi_V : in  std_logic_vector (7 downto 0);
    idata_176_roi_V : in  std_logic_vector (7 downto 0);
    idata_177_roi_V : in  std_logic_vector (7 downto 0);
    idata_178_roi_V : in  std_logic_vector (7 downto 0);
    idata_179_roi_V : in  std_logic_vector (7 downto 0);
    idata_180_roi_V : in  std_logic_vector (7 downto 0);
    idata_181_roi_V : in  std_logic_vector (7 downto 0);
    idata_182_roi_V : in  std_logic_vector (7 downto 0);
    idata_183_roi_V : in  std_logic_vector (7 downto 0);
    idata_184_roi_V : in  std_logic_vector (7 downto 0);
    idata_185_roi_V : in  std_logic_vector (7 downto 0);
    idata_186_roi_V : in  std_logic_vector (7 downto 0);
    idata_187_roi_V : in  std_logic_vector (7 downto 0);
    idata_188_roi_V : in  std_logic_vector (7 downto 0);
    idata_189_roi_V : in  std_logic_vector (7 downto 0);
    idata_190_roi_V : in  std_logic_vector (7 downto 0);
    idata_191_roi_V : in  std_logic_vector (7 downto 0);
    idata_192_roi_V : in  std_logic_vector (7 downto 0);
    idata_193_roi_V : in  std_logic_vector (7 downto 0);
    idata_194_roi_V : in  std_logic_vector (7 downto 0);
    idata_195_roi_V : in  std_logic_vector (7 downto 0);
    idata_196_roi_V : in  std_logic_vector (7 downto 0);
    idata_197_roi_V : in  std_logic_vector (7 downto 0);
    idata_198_roi_V : in  std_logic_vector (7 downto 0);
    idata_199_roi_V : in  std_logic_vector (7 downto 0);
    idata_200_roi_V : in  std_logic_vector (7 downto 0);
    idata_201_roi_V : in  std_logic_vector (7 downto 0);
    idata_202_roi_V : in  std_logic_vector (7 downto 0);
    idata_203_roi_V : in  std_logic_vector (7 downto 0);
    idata_204_roi_V : in  std_logic_vector (7 downto 0);
    idata_205_roi_V : in  std_logic_vector (7 downto 0);
    idata_206_roi_V : in  std_logic_vector (7 downto 0);
    idata_207_roi_V : in  std_logic_vector (7 downto 0);
    idata_208_roi_V : in  std_logic_vector (7 downto 0);
    idata_209_roi_V : in  std_logic_vector (7 downto 0);
    idata_210_roi_V : in  std_logic_vector (7 downto 0);
    idata_211_roi_V : in  std_logic_vector (7 downto 0);
    idata_212_roi_V : in  std_logic_vector (7 downto 0);
    idata_213_roi_V : in  std_logic_vector (7 downto 0);
    idata_214_roi_V : in  std_logic_vector (7 downto 0);
    idata_215_roi_V : in  std_logic_vector (7 downto 0);
    idata_216_roi_V : in  std_logic_vector (7 downto 0);
    idata_217_roi_V : in  std_logic_vector (7 downto 0);
    idata_218_roi_V : in  std_logic_vector (7 downto 0);
    idata_219_roi_V : in  std_logic_vector (7 downto 0);
    idata_220_roi_V : in  std_logic_vector (7 downto 0);
    idata_221_roi_V : in  std_logic_vector (7 downto 0);
    idata_222_roi_V : in  std_logic_vector (7 downto 0);
    idata_223_roi_V : in  std_logic_vector (7 downto 0);
    idata_224_roi_V : in  std_logic_vector (7 downto 0);
    idata_225_roi_V : in  std_logic_vector (7 downto 0);
    idata_226_roi_V : in  std_logic_vector (7 downto 0);
    idata_227_roi_V : in  std_logic_vector (7 downto 0);
    idata_228_roi_V : in  std_logic_vector (7 downto 0);
    idata_229_roi_V : in  std_logic_vector (7 downto 0);
    idata_230_roi_V : in  std_logic_vector (7 downto 0);
    idata_231_roi_V : in  std_logic_vector (7 downto 0);
    idata_232_roi_V : in  std_logic_vector (7 downto 0);
    idata_233_roi_V : in  std_logic_vector (7 downto 0);
    idata_234_roi_V : in  std_logic_vector (7 downto 0);
    idata_235_roi_V : in  std_logic_vector (7 downto 0);
    idata_236_roi_V : in  std_logic_vector (7 downto 0);
    idata_237_roi_V : in  std_logic_vector (7 downto 0);
    idata_238_roi_V : in  std_logic_vector (7 downto 0);
    idata_239_roi_V : in  std_logic_vector (7 downto 0);
    idata_240_roi_V : in  std_logic_vector (7 downto 0);
    idata_241_roi_V : in  std_logic_vector (7 downto 0);
    idata_242_roi_V : in  std_logic_vector (7 downto 0);
    idata_243_roi_V : in  std_logic_vector (7 downto 0);
    idata_244_roi_V : in  std_logic_vector (7 downto 0);
    idata_245_roi_V : in  std_logic_vector (7 downto 0);
    idata_246_roi_V : in  std_logic_vector (7 downto 0);
    idata_247_roi_V : in  std_logic_vector (7 downto 0);
    idata_248_roi_V : in  std_logic_vector (7 downto 0);
    idata_249_roi_V : in  std_logic_vector (7 downto 0);
    idata_250_roi_V : in  std_logic_vector (7 downto 0);
    idata_251_roi_V : in  std_logic_vector (7 downto 0);
    idata_252_roi_V : in  std_logic_vector (7 downto 0);
    idata_253_roi_V : in  std_logic_vector (7 downto 0);
    idata_254_roi_V : in  std_logic_vector (7 downto 0);
    idata_255_roi_V : in  std_logic_vector (7 downto 0);
    idata_256_roi_V : in  std_logic_vector (7 downto 0);
    idata_257_roi_V : in  std_logic_vector (7 downto 0);
    idata_258_roi_V : in  std_logic_vector (7 downto 0);
    idata_259_roi_V : in  std_logic_vector (7 downto 0);
    idata_260_roi_V : in  std_logic_vector (7 downto 0);
    idata_261_roi_V : in  std_logic_vector (7 downto 0);
    idata_262_roi_V : in  std_logic_vector (7 downto 0);
    idata_263_roi_V : in  std_logic_vector (7 downto 0);
    idata_264_roi_V : in  std_logic_vector (7 downto 0);
    idata_265_roi_V : in  std_logic_vector (7 downto 0);
    idata_266_roi_V : in  std_logic_vector (7 downto 0);
    idata_267_roi_V : in  std_logic_vector (7 downto 0);
    idata_268_roi_V : in  std_logic_vector (7 downto 0);
    idata_269_roi_V : in  std_logic_vector (7 downto 0);
    idata_270_roi_V : in  std_logic_vector (7 downto 0);
    idata_271_roi_V : in  std_logic_vector (7 downto 0);
    idata_272_roi_V : in  std_logic_vector (7 downto 0);
    idata_273_roi_V : in  std_logic_vector (7 downto 0);
    idata_274_roi_V : in  std_logic_vector (7 downto 0);
    idata_275_roi_V : in  std_logic_vector (7 downto 0);
    idata_276_roi_V : in  std_logic_vector (7 downto 0);
    idata_277_roi_V : in  std_logic_vector (7 downto 0);
    idata_278_roi_V : in  std_logic_vector (7 downto 0);
    idata_279_roi_V : in  std_logic_vector (7 downto 0);
    idata_280_roi_V : in  std_logic_vector (7 downto 0);
    idata_281_roi_V : in  std_logic_vector (7 downto 0);
    idata_282_roi_V : in  std_logic_vector (7 downto 0);
    idata_283_roi_V : in  std_logic_vector (7 downto 0);
    idata_284_roi_V : in  std_logic_vector (7 downto 0);
    idata_285_roi_V : in  std_logic_vector (7 downto 0);
    idata_286_roi_V : in  std_logic_vector (7 downto 0);
    idata_287_roi_V : in  std_logic_vector (7 downto 0);
    idata_288_roi_V : in  std_logic_vector (7 downto 0);
    idata_289_roi_V : in  std_logic_vector (7 downto 0);
    idata_290_roi_V : in  std_logic_vector (7 downto 0);
    idata_291_roi_V : in  std_logic_vector (7 downto 0);
    idata_292_roi_V : in  std_logic_vector (7 downto 0);
    idata_293_roi_V : in  std_logic_vector (7 downto 0);
    idata_294_roi_V : in  std_logic_vector (7 downto 0);
    idata_295_roi_V : in  std_logic_vector (7 downto 0);
    idata_296_roi_V : in  std_logic_vector (7 downto 0);
    idata_297_roi_V : in  std_logic_vector (7 downto 0);
    idata_298_roi_V : in  std_logic_vector (7 downto 0);
    idata_299_roi_V : in  std_logic_vector (7 downto 0);
    idata_300_roi_V : in  std_logic_vector (7 downto 0);
    idata_301_roi_V : in  std_logic_vector (7 downto 0);
    idata_302_roi_V : in  std_logic_vector (7 downto 0);
    idata_303_roi_V : in  std_logic_vector (7 downto 0);
    idata_304_roi_V : in  std_logic_vector (7 downto 0);
    idata_305_roi_V : in  std_logic_vector (7 downto 0);
    idata_306_roi_V : in  std_logic_vector (7 downto 0);
    idata_307_roi_V : in  std_logic_vector (7 downto 0);
    idata_308_roi_V : in  std_logic_vector (7 downto 0);
    idata_309_roi_V : in  std_logic_vector (7 downto 0);
    idata_310_roi_V : in  std_logic_vector (7 downto 0);
    idata_311_roi_V : in  std_logic_vector (7 downto 0);
    idata_312_roi_V : in  std_logic_vector (7 downto 0);
    idata_313_roi_V : in  std_logic_vector (7 downto 0);
    idata_314_roi_V : in  std_logic_vector (7 downto 0);
    idata_315_roi_V : in  std_logic_vector (7 downto 0);
    idata_316_roi_V : in  std_logic_vector (7 downto 0);
    idata_317_roi_V : in  std_logic_vector (7 downto 0);
    idata_318_roi_V : in  std_logic_vector (7 downto 0);
    idata_319_roi_V : in  std_logic_vector (7 downto 0);
    idata_320_roi_V : in  std_logic_vector (7 downto 0);
    idata_321_roi_V : in  std_logic_vector (7 downto 0);
    idata_322_roi_V : in  std_logic_vector (7 downto 0);
    idata_323_roi_V : in  std_logic_vector (7 downto 0);
    idata_324_roi_V : in  std_logic_vector (7 downto 0);
    idata_325_roi_V : in  std_logic_vector (7 downto 0);
    idata_326_roi_V : in  std_logic_vector (7 downto 0);
    idata_327_roi_V : in  std_logic_vector (7 downto 0);
    idata_328_roi_V : in  std_logic_vector (7 downto 0);
    idata_329_roi_V : in  std_logic_vector (7 downto 0);
    idata_330_roi_V : in  std_logic_vector (7 downto 0);
    idata_331_roi_V : in  std_logic_vector (7 downto 0);
    idata_332_roi_V : in  std_logic_vector (7 downto 0);
    idata_333_roi_V : in  std_logic_vector (7 downto 0);
    idata_334_roi_V : in  std_logic_vector (7 downto 0);
    idata_335_roi_V : in  std_logic_vector (7 downto 0);
    idata_336_roi_V : in  std_logic_vector (7 downto 0);
    idata_337_roi_V : in  std_logic_vector (7 downto 0);
    idata_338_roi_V : in  std_logic_vector (7 downto 0);
    idata_339_roi_V : in  std_logic_vector (7 downto 0);
    idata_340_roi_V : in  std_logic_vector (7 downto 0);
    idata_341_roi_V : in  std_logic_vector (7 downto 0);
    idata_342_roi_V : in  std_logic_vector (7 downto 0);
    idata_343_roi_V : in  std_logic_vector (7 downto 0);
    idata_344_roi_V : in  std_logic_vector (7 downto 0);
    idata_345_roi_V : in  std_logic_vector (7 downto 0);
    idata_346_roi_V : in  std_logic_vector (7 downto 0);
    idata_347_roi_V : in  std_logic_vector (7 downto 0);
    idata_348_roi_V : in  std_logic_vector (7 downto 0);
    idata_349_roi_V : in  std_logic_vector (7 downto 0);
    idata_350_roi_V : in  std_logic_vector (7 downto 0);
    idata_351_roi_V : in  std_logic_vector (7 downto 0);
    idata_0_flg_V   : in  std_logic_vector (3 downto 0);
    idata_1_flg_V   : in  std_logic_vector (3 downto 0);
    idata_2_flg_V   : in  std_logic_vector (3 downto 0);
    idata_3_flg_V   : in  std_logic_vector (3 downto 0);
    idata_4_flg_V   : in  std_logic_vector (3 downto 0);
    idata_5_flg_V   : in  std_logic_vector (3 downto 0);
    idata_6_flg_V   : in  std_logic_vector (3 downto 0);
    idata_7_flg_V   : in  std_logic_vector (3 downto 0);
    idata_8_flg_V   : in  std_logic_vector (3 downto 0);
    idata_9_flg_V   : in  std_logic_vector (3 downto 0);
    idata_10_flg_V  : in  std_logic_vector (3 downto 0);
    idata_11_flg_V  : in  std_logic_vector (3 downto 0);
    idata_12_flg_V  : in  std_logic_vector (3 downto 0);
    idata_13_flg_V  : in  std_logic_vector (3 downto 0);
    idata_14_flg_V  : in  std_logic_vector (3 downto 0);
    idata_15_flg_V  : in  std_logic_vector (3 downto 0);
    idata_16_flg_V  : in  std_logic_vector (3 downto 0);
    idata_17_flg_V  : in  std_logic_vector (3 downto 0);
    idata_18_flg_V  : in  std_logic_vector (3 downto 0);
    idata_19_flg_V  : in  std_logic_vector (3 downto 0);
    idata_20_flg_V  : in  std_logic_vector (3 downto 0);
    idata_21_flg_V  : in  std_logic_vector (3 downto 0);
    idata_22_flg_V  : in  std_logic_vector (3 downto 0);
    idata_23_flg_V  : in  std_logic_vector (3 downto 0);
    idata_24_flg_V  : in  std_logic_vector (3 downto 0);
    idata_25_flg_V  : in  std_logic_vector (3 downto 0);
    idata_26_flg_V  : in  std_logic_vector (3 downto 0);
    idata_27_flg_V  : in  std_logic_vector (3 downto 0);
    idata_28_flg_V  : in  std_logic_vector (3 downto 0);
    idata_29_flg_V  : in  std_logic_vector (3 downto 0);
    idata_30_flg_V  : in  std_logic_vector (3 downto 0);
    idata_31_flg_V  : in  std_logic_vector (3 downto 0);
    idata_32_flg_V  : in  std_logic_vector (3 downto 0);
    idata_33_flg_V  : in  std_logic_vector (3 downto 0);
    idata_34_flg_V  : in  std_logic_vector (3 downto 0);
    idata_35_flg_V  : in  std_logic_vector (3 downto 0);
    idata_36_flg_V  : in  std_logic_vector (3 downto 0);
    idata_37_flg_V  : in  std_logic_vector (3 downto 0);
    idata_38_flg_V  : in  std_logic_vector (3 downto 0);
    idata_39_flg_V  : in  std_logic_vector (3 downto 0);
    idata_40_flg_V  : in  std_logic_vector (3 downto 0);
    idata_41_flg_V  : in  std_logic_vector (3 downto 0);
    idata_42_flg_V  : in  std_logic_vector (3 downto 0);
    idata_43_flg_V  : in  std_logic_vector (3 downto 0);
    idata_44_flg_V  : in  std_logic_vector (3 downto 0);
    idata_45_flg_V  : in  std_logic_vector (3 downto 0);
    idata_46_flg_V  : in  std_logic_vector (3 downto 0);
    idata_47_flg_V  : in  std_logic_vector (3 downto 0);
    idata_48_flg_V  : in  std_logic_vector (3 downto 0);
    idata_49_flg_V  : in  std_logic_vector (3 downto 0);
    idata_50_flg_V  : in  std_logic_vector (3 downto 0);
    idata_51_flg_V  : in  std_logic_vector (3 downto 0);
    idata_52_flg_V  : in  std_logic_vector (3 downto 0);
    idata_53_flg_V  : in  std_logic_vector (3 downto 0);
    idata_54_flg_V  : in  std_logic_vector (3 downto 0);
    idata_55_flg_V  : in  std_logic_vector (3 downto 0);
    idata_56_flg_V  : in  std_logic_vector (3 downto 0);
    idata_57_flg_V  : in  std_logic_vector (3 downto 0);
    idata_58_flg_V  : in  std_logic_vector (3 downto 0);
    idata_59_flg_V  : in  std_logic_vector (3 downto 0);
    idata_60_flg_V  : in  std_logic_vector (3 downto 0);
    idata_61_flg_V  : in  std_logic_vector (3 downto 0);
    idata_62_flg_V  : in  std_logic_vector (3 downto 0);
    idata_63_flg_V  : in  std_logic_vector (3 downto 0);
    idata_64_flg_V  : in  std_logic_vector (3 downto 0);
    idata_65_flg_V  : in  std_logic_vector (3 downto 0);
    idata_66_flg_V  : in  std_logic_vector (3 downto 0);
    idata_67_flg_V  : in  std_logic_vector (3 downto 0);
    idata_68_flg_V  : in  std_logic_vector (3 downto 0);
    idata_69_flg_V  : in  std_logic_vector (3 downto 0);
    idata_70_flg_V  : in  std_logic_vector (3 downto 0);
    idata_71_flg_V  : in  std_logic_vector (3 downto 0);
    idata_72_flg_V  : in  std_logic_vector (3 downto 0);
    idata_73_flg_V  : in  std_logic_vector (3 downto 0);
    idata_74_flg_V  : in  std_logic_vector (3 downto 0);
    idata_75_flg_V  : in  std_logic_vector (3 downto 0);
    idata_76_flg_V  : in  std_logic_vector (3 downto 0);
    idata_77_flg_V  : in  std_logic_vector (3 downto 0);
    idata_78_flg_V  : in  std_logic_vector (3 downto 0);
    idata_79_flg_V  : in  std_logic_vector (3 downto 0);
    idata_80_flg_V  : in  std_logic_vector (3 downto 0);
    idata_81_flg_V  : in  std_logic_vector (3 downto 0);
    idata_82_flg_V  : in  std_logic_vector (3 downto 0);
    idata_83_flg_V  : in  std_logic_vector (3 downto 0);
    idata_84_flg_V  : in  std_logic_vector (3 downto 0);
    idata_85_flg_V  : in  std_logic_vector (3 downto 0);
    idata_86_flg_V  : in  std_logic_vector (3 downto 0);
    idata_87_flg_V  : in  std_logic_vector (3 downto 0);
    idata_88_flg_V  : in  std_logic_vector (3 downto 0);
    idata_89_flg_V  : in  std_logic_vector (3 downto 0);
    idata_90_flg_V  : in  std_logic_vector (3 downto 0);
    idata_91_flg_V  : in  std_logic_vector (3 downto 0);
    idata_92_flg_V  : in  std_logic_vector (3 downto 0);
    idata_93_flg_V  : in  std_logic_vector (3 downto 0);
    idata_94_flg_V  : in  std_logic_vector (3 downto 0);
    idata_95_flg_V  : in  std_logic_vector (3 downto 0);
    idata_96_flg_V  : in  std_logic_vector (3 downto 0);
    idata_97_flg_V  : in  std_logic_vector (3 downto 0);
    idata_98_flg_V  : in  std_logic_vector (3 downto 0);
    idata_99_flg_V  : in  std_logic_vector (3 downto 0);
    idata_100_flg_V : in  std_logic_vector (3 downto 0);
    idata_101_flg_V : in  std_logic_vector (3 downto 0);
    idata_102_flg_V : in  std_logic_vector (3 downto 0);
    idata_103_flg_V : in  std_logic_vector (3 downto 0);
    idata_104_flg_V : in  std_logic_vector (3 downto 0);
    idata_105_flg_V : in  std_logic_vector (3 downto 0);
    idata_106_flg_V : in  std_logic_vector (3 downto 0);
    idata_107_flg_V : in  std_logic_vector (3 downto 0);
    idata_108_flg_V : in  std_logic_vector (3 downto 0);
    idata_109_flg_V : in  std_logic_vector (3 downto 0);
    idata_110_flg_V : in  std_logic_vector (3 downto 0);
    idata_111_flg_V : in  std_logic_vector (3 downto 0);
    idata_112_flg_V : in  std_logic_vector (3 downto 0);
    idata_113_flg_V : in  std_logic_vector (3 downto 0);
    idata_114_flg_V : in  std_logic_vector (3 downto 0);
    idata_115_flg_V : in  std_logic_vector (3 downto 0);
    idata_116_flg_V : in  std_logic_vector (3 downto 0);
    idata_117_flg_V : in  std_logic_vector (3 downto 0);
    idata_118_flg_V : in  std_logic_vector (3 downto 0);
    idata_119_flg_V : in  std_logic_vector (3 downto 0);
    idata_120_flg_V : in  std_logic_vector (3 downto 0);
    idata_121_flg_V : in  std_logic_vector (3 downto 0);
    idata_122_flg_V : in  std_logic_vector (3 downto 0);
    idata_123_flg_V : in  std_logic_vector (3 downto 0);
    idata_124_flg_V : in  std_logic_vector (3 downto 0);
    idata_125_flg_V : in  std_logic_vector (3 downto 0);
    idata_126_flg_V : in  std_logic_vector (3 downto 0);
    idata_127_flg_V : in  std_logic_vector (3 downto 0);
    idata_128_flg_V : in  std_logic_vector (3 downto 0);
    idata_129_flg_V : in  std_logic_vector (3 downto 0);
    idata_130_flg_V : in  std_logic_vector (3 downto 0);
    idata_131_flg_V : in  std_logic_vector (3 downto 0);
    idata_132_flg_V : in  std_logic_vector (3 downto 0);
    idata_133_flg_V : in  std_logic_vector (3 downto 0);
    idata_134_flg_V : in  std_logic_vector (3 downto 0);
    idata_135_flg_V : in  std_logic_vector (3 downto 0);
    idata_136_flg_V : in  std_logic_vector (3 downto 0);
    idata_137_flg_V : in  std_logic_vector (3 downto 0);
    idata_138_flg_V : in  std_logic_vector (3 downto 0);
    idata_139_flg_V : in  std_logic_vector (3 downto 0);
    idata_140_flg_V : in  std_logic_vector (3 downto 0);
    idata_141_flg_V : in  std_logic_vector (3 downto 0);
    idata_142_flg_V : in  std_logic_vector (3 downto 0);
    idata_143_flg_V : in  std_logic_vector (3 downto 0);
    idata_144_flg_V : in  std_logic_vector (3 downto 0);
    idata_145_flg_V : in  std_logic_vector (3 downto 0);
    idata_146_flg_V : in  std_logic_vector (3 downto 0);
    idata_147_flg_V : in  std_logic_vector (3 downto 0);
    idata_148_flg_V : in  std_logic_vector (3 downto 0);
    idata_149_flg_V : in  std_logic_vector (3 downto 0);
    idata_150_flg_V : in  std_logic_vector (3 downto 0);
    idata_151_flg_V : in  std_logic_vector (3 downto 0);
    idata_152_flg_V : in  std_logic_vector (3 downto 0);
    idata_153_flg_V : in  std_logic_vector (3 downto 0);
    idata_154_flg_V : in  std_logic_vector (3 downto 0);
    idata_155_flg_V : in  std_logic_vector (3 downto 0);
    idata_156_flg_V : in  std_logic_vector (3 downto 0);
    idata_157_flg_V : in  std_logic_vector (3 downto 0);
    idata_158_flg_V : in  std_logic_vector (3 downto 0);
    idata_159_flg_V : in  std_logic_vector (3 downto 0);
    idata_160_flg_V : in  std_logic_vector (3 downto 0);
    idata_161_flg_V : in  std_logic_vector (3 downto 0);
    idata_162_flg_V : in  std_logic_vector (3 downto 0);
    idata_163_flg_V : in  std_logic_vector (3 downto 0);
    idata_164_flg_V : in  std_logic_vector (3 downto 0);
    idata_165_flg_V : in  std_logic_vector (3 downto 0);
    idata_166_flg_V : in  std_logic_vector (3 downto 0);
    idata_167_flg_V : in  std_logic_vector (3 downto 0);
    idata_168_flg_V : in  std_logic_vector (3 downto 0);
    idata_169_flg_V : in  std_logic_vector (3 downto 0);
    idata_170_flg_V : in  std_logic_vector (3 downto 0);
    idata_171_flg_V : in  std_logic_vector (3 downto 0);
    idata_172_flg_V : in  std_logic_vector (3 downto 0);
    idata_173_flg_V : in  std_logic_vector (3 downto 0);
    idata_174_flg_V : in  std_logic_vector (3 downto 0);
    idata_175_flg_V : in  std_logic_vector (3 downto 0);
    idata_176_flg_V : in  std_logic_vector (3 downto 0);
    idata_177_flg_V : in  std_logic_vector (3 downto 0);
    idata_178_flg_V : in  std_logic_vector (3 downto 0);
    idata_179_flg_V : in  std_logic_vector (3 downto 0);
    idata_180_flg_V : in  std_logic_vector (3 downto 0);
    idata_181_flg_V : in  std_logic_vector (3 downto 0);
    idata_182_flg_V : in  std_logic_vector (3 downto 0);
    idata_183_flg_V : in  std_logic_vector (3 downto 0);
    idata_184_flg_V : in  std_logic_vector (3 downto 0);
    idata_185_flg_V : in  std_logic_vector (3 downto 0);
    idata_186_flg_V : in  std_logic_vector (3 downto 0);
    idata_187_flg_V : in  std_logic_vector (3 downto 0);
    idata_188_flg_V : in  std_logic_vector (3 downto 0);
    idata_189_flg_V : in  std_logic_vector (3 downto 0);
    idata_190_flg_V : in  std_logic_vector (3 downto 0);
    idata_191_flg_V : in  std_logic_vector (3 downto 0);
    idata_192_flg_V : in  std_logic_vector (3 downto 0);
    idata_193_flg_V : in  std_logic_vector (3 downto 0);
    idata_194_flg_V : in  std_logic_vector (3 downto 0);
    idata_195_flg_V : in  std_logic_vector (3 downto 0);
    idata_196_flg_V : in  std_logic_vector (3 downto 0);
    idata_197_flg_V : in  std_logic_vector (3 downto 0);
    idata_198_flg_V : in  std_logic_vector (3 downto 0);
    idata_199_flg_V : in  std_logic_vector (3 downto 0);
    idata_200_flg_V : in  std_logic_vector (3 downto 0);
    idata_201_flg_V : in  std_logic_vector (3 downto 0);
    idata_202_flg_V : in  std_logic_vector (3 downto 0);
    idata_203_flg_V : in  std_logic_vector (3 downto 0);
    idata_204_flg_V : in  std_logic_vector (3 downto 0);
    idata_205_flg_V : in  std_logic_vector (3 downto 0);
    idata_206_flg_V : in  std_logic_vector (3 downto 0);
    idata_207_flg_V : in  std_logic_vector (3 downto 0);
    idata_208_flg_V : in  std_logic_vector (3 downto 0);
    idata_209_flg_V : in  std_logic_vector (3 downto 0);
    idata_210_flg_V : in  std_logic_vector (3 downto 0);
    idata_211_flg_V : in  std_logic_vector (3 downto 0);
    idata_212_flg_V : in  std_logic_vector (3 downto 0);
    idata_213_flg_V : in  std_logic_vector (3 downto 0);
    idata_214_flg_V : in  std_logic_vector (3 downto 0);
    idata_215_flg_V : in  std_logic_vector (3 downto 0);
    idata_216_flg_V : in  std_logic_vector (3 downto 0);
    idata_217_flg_V : in  std_logic_vector (3 downto 0);
    idata_218_flg_V : in  std_logic_vector (3 downto 0);
    idata_219_flg_V : in  std_logic_vector (3 downto 0);
    idata_220_flg_V : in  std_logic_vector (3 downto 0);
    idata_221_flg_V : in  std_logic_vector (3 downto 0);
    idata_222_flg_V : in  std_logic_vector (3 downto 0);
    idata_223_flg_V : in  std_logic_vector (3 downto 0);
    idata_224_flg_V : in  std_logic_vector (3 downto 0);
    idata_225_flg_V : in  std_logic_vector (3 downto 0);
    idata_226_flg_V : in  std_logic_vector (3 downto 0);
    idata_227_flg_V : in  std_logic_vector (3 downto 0);
    idata_228_flg_V : in  std_logic_vector (3 downto 0);
    idata_229_flg_V : in  std_logic_vector (3 downto 0);
    idata_230_flg_V : in  std_logic_vector (3 downto 0);
    idata_231_flg_V : in  std_logic_vector (3 downto 0);
    idata_232_flg_V : in  std_logic_vector (3 downto 0);
    idata_233_flg_V : in  std_logic_vector (3 downto 0);
    idata_234_flg_V : in  std_logic_vector (3 downto 0);
    idata_235_flg_V : in  std_logic_vector (3 downto 0);
    idata_236_flg_V : in  std_logic_vector (3 downto 0);
    idata_237_flg_V : in  std_logic_vector (3 downto 0);
    idata_238_flg_V : in  std_logic_vector (3 downto 0);
    idata_239_flg_V : in  std_logic_vector (3 downto 0);
    idata_240_flg_V : in  std_logic_vector (3 downto 0);
    idata_241_flg_V : in  std_logic_vector (3 downto 0);
    idata_242_flg_V : in  std_logic_vector (3 downto 0);
    idata_243_flg_V : in  std_logic_vector (3 downto 0);
    idata_244_flg_V : in  std_logic_vector (3 downto 0);
    idata_245_flg_V : in  std_logic_vector (3 downto 0);
    idata_246_flg_V : in  std_logic_vector (3 downto 0);
    idata_247_flg_V : in  std_logic_vector (3 downto 0);
    idata_248_flg_V : in  std_logic_vector (3 downto 0);
    idata_249_flg_V : in  std_logic_vector (3 downto 0);
    idata_250_flg_V : in  std_logic_vector (3 downto 0);
    idata_251_flg_V : in  std_logic_vector (3 downto 0);
    idata_252_flg_V : in  std_logic_vector (3 downto 0);
    idata_253_flg_V : in  std_logic_vector (3 downto 0);
    idata_254_flg_V : in  std_logic_vector (3 downto 0);
    idata_255_flg_V : in  std_logic_vector (3 downto 0);
    idata_256_flg_V : in  std_logic_vector (3 downto 0);
    idata_257_flg_V : in  std_logic_vector (3 downto 0);
    idata_258_flg_V : in  std_logic_vector (3 downto 0);
    idata_259_flg_V : in  std_logic_vector (3 downto 0);
    idata_260_flg_V : in  std_logic_vector (3 downto 0);
    idata_261_flg_V : in  std_logic_vector (3 downto 0);
    idata_262_flg_V : in  std_logic_vector (3 downto 0);
    idata_263_flg_V : in  std_logic_vector (3 downto 0);
    idata_264_flg_V : in  std_logic_vector (3 downto 0);
    idata_265_flg_V : in  std_logic_vector (3 downto 0);
    idata_266_flg_V : in  std_logic_vector (3 downto 0);
    idata_267_flg_V : in  std_logic_vector (3 downto 0);
    idata_268_flg_V : in  std_logic_vector (3 downto 0);
    idata_269_flg_V : in  std_logic_vector (3 downto 0);
    idata_270_flg_V : in  std_logic_vector (3 downto 0);
    idata_271_flg_V : in  std_logic_vector (3 downto 0);
    idata_272_flg_V : in  std_logic_vector (3 downto 0);
    idata_273_flg_V : in  std_logic_vector (3 downto 0);
    idata_274_flg_V : in  std_logic_vector (3 downto 0);
    idata_275_flg_V : in  std_logic_vector (3 downto 0);
    idata_276_flg_V : in  std_logic_vector (3 downto 0);
    idata_277_flg_V : in  std_logic_vector (3 downto 0);
    idata_278_flg_V : in  std_logic_vector (3 downto 0);
    idata_279_flg_V : in  std_logic_vector (3 downto 0);
    idata_280_flg_V : in  std_logic_vector (3 downto 0);
    idata_281_flg_V : in  std_logic_vector (3 downto 0);
    idata_282_flg_V : in  std_logic_vector (3 downto 0);
    idata_283_flg_V : in  std_logic_vector (3 downto 0);
    idata_284_flg_V : in  std_logic_vector (3 downto 0);
    idata_285_flg_V : in  std_logic_vector (3 downto 0);
    idata_286_flg_V : in  std_logic_vector (3 downto 0);
    idata_287_flg_V : in  std_logic_vector (3 downto 0);
    idata_288_flg_V : in  std_logic_vector (3 downto 0);
    idata_289_flg_V : in  std_logic_vector (3 downto 0);
    idata_290_flg_V : in  std_logic_vector (3 downto 0);
    idata_291_flg_V : in  std_logic_vector (3 downto 0);
    idata_292_flg_V : in  std_logic_vector (3 downto 0);
    idata_293_flg_V : in  std_logic_vector (3 downto 0);
    idata_294_flg_V : in  std_logic_vector (3 downto 0);
    idata_295_flg_V : in  std_logic_vector (3 downto 0);
    idata_296_flg_V : in  std_logic_vector (3 downto 0);
    idata_297_flg_V : in  std_logic_vector (3 downto 0);
    idata_298_flg_V : in  std_logic_vector (3 downto 0);
    idata_299_flg_V : in  std_logic_vector (3 downto 0);
    idata_300_flg_V : in  std_logic_vector (3 downto 0);
    idata_301_flg_V : in  std_logic_vector (3 downto 0);
    idata_302_flg_V : in  std_logic_vector (3 downto 0);
    idata_303_flg_V : in  std_logic_vector (3 downto 0);
    idata_304_flg_V : in  std_logic_vector (3 downto 0);
    idata_305_flg_V : in  std_logic_vector (3 downto 0);
    idata_306_flg_V : in  std_logic_vector (3 downto 0);
    idata_307_flg_V : in  std_logic_vector (3 downto 0);
    idata_308_flg_V : in  std_logic_vector (3 downto 0);
    idata_309_flg_V : in  std_logic_vector (3 downto 0);
    idata_310_flg_V : in  std_logic_vector (3 downto 0);
    idata_311_flg_V : in  std_logic_vector (3 downto 0);
    idata_312_flg_V : in  std_logic_vector (3 downto 0);
    idata_313_flg_V : in  std_logic_vector (3 downto 0);
    idata_314_flg_V : in  std_logic_vector (3 downto 0);
    idata_315_flg_V : in  std_logic_vector (3 downto 0);
    idata_316_flg_V : in  std_logic_vector (3 downto 0);
    idata_317_flg_V : in  std_logic_vector (3 downto 0);
    idata_318_flg_V : in  std_logic_vector (3 downto 0);
    idata_319_flg_V : in  std_logic_vector (3 downto 0);
    idata_320_flg_V : in  std_logic_vector (3 downto 0);
    idata_321_flg_V : in  std_logic_vector (3 downto 0);
    idata_322_flg_V : in  std_logic_vector (3 downto 0);
    idata_323_flg_V : in  std_logic_vector (3 downto 0);
    idata_324_flg_V : in  std_logic_vector (3 downto 0);
    idata_325_flg_V : in  std_logic_vector (3 downto 0);
    idata_326_flg_V : in  std_logic_vector (3 downto 0);
    idata_327_flg_V : in  std_logic_vector (3 downto 0);
    idata_328_flg_V : in  std_logic_vector (3 downto 0);
    idata_329_flg_V : in  std_logic_vector (3 downto 0);
    idata_330_flg_V : in  std_logic_vector (3 downto 0);
    idata_331_flg_V : in  std_logic_vector (3 downto 0);
    idata_332_flg_V : in  std_logic_vector (3 downto 0);
    idata_333_flg_V : in  std_logic_vector (3 downto 0);
    idata_334_flg_V : in  std_logic_vector (3 downto 0);
    idata_335_flg_V : in  std_logic_vector (3 downto 0);
    idata_336_flg_V : in  std_logic_vector (3 downto 0);
    idata_337_flg_V : in  std_logic_vector (3 downto 0);
    idata_338_flg_V : in  std_logic_vector (3 downto 0);
    idata_339_flg_V : in  std_logic_vector (3 downto 0);
    idata_340_flg_V : in  std_logic_vector (3 downto 0);
    idata_341_flg_V : in  std_logic_vector (3 downto 0);
    idata_342_flg_V : in  std_logic_vector (3 downto 0);
    idata_343_flg_V : in  std_logic_vector (3 downto 0);
    idata_344_flg_V : in  std_logic_vector (3 downto 0);
    idata_345_flg_V : in  std_logic_vector (3 downto 0);
    idata_346_flg_V : in  std_logic_vector (3 downto 0);
    idata_347_flg_V : in  std_logic_vector (3 downto 0);
    idata_348_flg_V : in  std_logic_vector (3 downto 0);
    idata_349_flg_V : in  std_logic_vector (3 downto 0);
    idata_350_flg_V : in  std_logic_vector (3 downto 0);
    idata_351_flg_V : in  std_logic_vector (3 downto 0);
    odata_0_id_V    : out std_logic_vector (8 downto 0);
    odata_1_id_V    : out std_logic_vector (8 downto 0);
    odata_2_id_V    : out std_logic_vector (8 downto 0);
    odata_3_id_V    : out std_logic_vector (8 downto 0);
    odata_4_id_V    : out std_logic_vector (8 downto 0);
    odata_5_id_V    : out std_logic_vector (8 downto 0);
    odata_6_id_V    : out std_logic_vector (8 downto 0);
    odata_7_id_V    : out std_logic_vector (8 downto 0);
    odata_8_id_V    : out std_logic_vector (8 downto 0);
    odata_9_id_V    : out std_logic_vector (8 downto 0);
    odata_10_id_V   : out std_logic_vector (8 downto 0);
    odata_11_id_V   : out std_logic_vector (8 downto 0);
    odata_12_id_V   : out std_logic_vector (8 downto 0);
    odata_13_id_V   : out std_logic_vector (8 downto 0);
    odata_14_id_V   : out std_logic_vector (8 downto 0);
    odata_15_id_V   : out std_logic_vector (8 downto 0);
    odata_0_pt_V    : out std_logic_vector (3 downto 0);
    odata_1_pt_V    : out std_logic_vector (3 downto 0);
    odata_2_pt_V    : out std_logic_vector (3 downto 0);
    odata_3_pt_V    : out std_logic_vector (3 downto 0);
    odata_4_pt_V    : out std_logic_vector (3 downto 0);
    odata_5_pt_V    : out std_logic_vector (3 downto 0);
    odata_6_pt_V    : out std_logic_vector (3 downto 0);
    odata_7_pt_V    : out std_logic_vector (3 downto 0);
    odata_8_pt_V    : out std_logic_vector (3 downto 0);
    odata_9_pt_V    : out std_logic_vector (3 downto 0);
    odata_10_pt_V   : out std_logic_vector (3 downto 0);
    odata_11_pt_V   : out std_logic_vector (3 downto 0);
    odata_12_pt_V   : out std_logic_vector (3 downto 0);
    odata_13_pt_V   : out std_logic_vector (3 downto 0);
    odata_14_pt_V   : out std_logic_vector (3 downto 0);
    odata_15_pt_V   : out std_logic_vector (3 downto 0);
    odata_0_roi_V   : out std_logic_vector (7 downto 0);
    odata_1_roi_V   : out std_logic_vector (7 downto 0);
    odata_2_roi_V   : out std_logic_vector (7 downto 0);
    odata_3_roi_V   : out std_logic_vector (7 downto 0);
    odata_4_roi_V   : out std_logic_vector (7 downto 0);
    odata_5_roi_V   : out std_logic_vector (7 downto 0);
    odata_6_roi_V   : out std_logic_vector (7 downto 0);
    odata_7_roi_V   : out std_logic_vector (7 downto 0);
    odata_8_roi_V   : out std_logic_vector (7 downto 0);
    odata_9_roi_V   : out std_logic_vector (7 downto 0);
    odata_10_roi_V  : out std_logic_vector (7 downto 0);
    odata_11_roi_V  : out std_logic_vector (7 downto 0);
    odata_12_roi_V  : out std_logic_vector (7 downto 0);
    odata_13_roi_V  : out std_logic_vector (7 downto 0);
    odata_14_roi_V  : out std_logic_vector (7 downto 0);
    odata_15_roi_V  : out std_logic_vector (7 downto 0);
    odata_0_flg_V   : out std_logic_vector (3 downto 0);
    odata_1_flg_V   : out std_logic_vector (3 downto 0);
    odata_2_flg_V   : out std_logic_vector (3 downto 0);
    odata_3_flg_V   : out std_logic_vector (3 downto 0);
    odata_4_flg_V   : out std_logic_vector (3 downto 0);
    odata_5_flg_V   : out std_logic_vector (3 downto 0);
    odata_6_flg_V   : out std_logic_vector (3 downto 0);
    odata_7_flg_V   : out std_logic_vector (3 downto 0);
    odata_8_flg_V   : out std_logic_vector (3 downto 0);
    odata_9_flg_V   : out std_logic_vector (3 downto 0);
    odata_10_flg_V  : out std_logic_vector (3 downto 0);
    odata_11_flg_V  : out std_logic_vector (3 downto 0);
    odata_12_flg_V  : out std_logic_vector (3 downto 0);
    odata_13_flg_V  : out std_logic_vector (3 downto 0);
    odata_14_flg_V  : out std_logic_vector (3 downto 0);
    odata_15_flg_V  : out std_logic_vector (3 downto 0));

end entity compare_wrapper;

architecture rtl of compare_wrapper is

  component compare_main is
    port (
      ap_clk          : in  std_logic;
      ap_rst          : in  std_logic;
      ap_start        : in  std_logic;
      ap_done         : out std_logic;
      ap_idle         : out std_logic;
      ap_ready        : out std_logic;
      idata_0_pt_V    : in  std_logic_vector (3 downto 0);
      idata_1_pt_V    : in  std_logic_vector (3 downto 0);
      idata_2_pt_V    : in  std_logic_vector (3 downto 0);
      idata_3_pt_V    : in  std_logic_vector (3 downto 0);
      idata_4_pt_V    : in  std_logic_vector (3 downto 0);
      idata_5_pt_V    : in  std_logic_vector (3 downto 0);
      idata_6_pt_V    : in  std_logic_vector (3 downto 0);
      idata_7_pt_V    : in  std_logic_vector (3 downto 0);
      idata_8_pt_V    : in  std_logic_vector (3 downto 0);
      idata_9_pt_V    : in  std_logic_vector (3 downto 0);
      idata_10_pt_V   : in  std_logic_vector (3 downto 0);
      idata_11_pt_V   : in  std_logic_vector (3 downto 0);
      idata_12_pt_V   : in  std_logic_vector (3 downto 0);
      idata_13_pt_V   : in  std_logic_vector (3 downto 0);
      idata_14_pt_V   : in  std_logic_vector (3 downto 0);
      idata_15_pt_V   : in  std_logic_vector (3 downto 0);
      idata_16_pt_V   : in  std_logic_vector (3 downto 0);
      idata_17_pt_V   : in  std_logic_vector (3 downto 0);
      idata_18_pt_V   : in  std_logic_vector (3 downto 0);
      idata_19_pt_V   : in  std_logic_vector (3 downto 0);
      idata_20_pt_V   : in  std_logic_vector (3 downto 0);
      idata_21_pt_V   : in  std_logic_vector (3 downto 0);
      idata_22_pt_V   : in  std_logic_vector (3 downto 0);
      idata_23_pt_V   : in  std_logic_vector (3 downto 0);
      idata_24_pt_V   : in  std_logic_vector (3 downto 0);
      idata_25_pt_V   : in  std_logic_vector (3 downto 0);
      idata_26_pt_V   : in  std_logic_vector (3 downto 0);
      idata_27_pt_V   : in  std_logic_vector (3 downto 0);
      idata_28_pt_V   : in  std_logic_vector (3 downto 0);
      idata_29_pt_V   : in  std_logic_vector (3 downto 0);
      idata_30_pt_V   : in  std_logic_vector (3 downto 0);
      idata_31_pt_V   : in  std_logic_vector (3 downto 0);
      idata_32_pt_V   : in  std_logic_vector (3 downto 0);
      idata_33_pt_V   : in  std_logic_vector (3 downto 0);
      idata_34_pt_V   : in  std_logic_vector (3 downto 0);
      idata_35_pt_V   : in  std_logic_vector (3 downto 0);
      idata_36_pt_V   : in  std_logic_vector (3 downto 0);
      idata_37_pt_V   : in  std_logic_vector (3 downto 0);
      idata_38_pt_V   : in  std_logic_vector (3 downto 0);
      idata_39_pt_V   : in  std_logic_vector (3 downto 0);
      idata_40_pt_V   : in  std_logic_vector (3 downto 0);
      idata_41_pt_V   : in  std_logic_vector (3 downto 0);
      idata_42_pt_V   : in  std_logic_vector (3 downto 0);
      idata_43_pt_V   : in  std_logic_vector (3 downto 0);
      idata_44_pt_V   : in  std_logic_vector (3 downto 0);
      idata_45_pt_V   : in  std_logic_vector (3 downto 0);
      idata_46_pt_V   : in  std_logic_vector (3 downto 0);
      idata_47_pt_V   : in  std_logic_vector (3 downto 0);
      idata_48_pt_V   : in  std_logic_vector (3 downto 0);
      idata_49_pt_V   : in  std_logic_vector (3 downto 0);
      idata_50_pt_V   : in  std_logic_vector (3 downto 0);
      idata_51_pt_V   : in  std_logic_vector (3 downto 0);
      idata_52_pt_V   : in  std_logic_vector (3 downto 0);
      idata_53_pt_V   : in  std_logic_vector (3 downto 0);
      idata_54_pt_V   : in  std_logic_vector (3 downto 0);
      idata_55_pt_V   : in  std_logic_vector (3 downto 0);
      idata_56_pt_V   : in  std_logic_vector (3 downto 0);
      idata_57_pt_V   : in  std_logic_vector (3 downto 0);
      idata_58_pt_V   : in  std_logic_vector (3 downto 0);
      idata_59_pt_V   : in  std_logic_vector (3 downto 0);
      idata_60_pt_V   : in  std_logic_vector (3 downto 0);
      idata_61_pt_V   : in  std_logic_vector (3 downto 0);
      idata_62_pt_V   : in  std_logic_vector (3 downto 0);
      idata_63_pt_V   : in  std_logic_vector (3 downto 0);
      idata_64_pt_V   : in  std_logic_vector (3 downto 0);
      idata_65_pt_V   : in  std_logic_vector (3 downto 0);
      idata_66_pt_V   : in  std_logic_vector (3 downto 0);
      idata_67_pt_V   : in  std_logic_vector (3 downto 0);
      idata_68_pt_V   : in  std_logic_vector (3 downto 0);
      idata_69_pt_V   : in  std_logic_vector (3 downto 0);
      idata_70_pt_V   : in  std_logic_vector (3 downto 0);
      idata_71_pt_V   : in  std_logic_vector (3 downto 0);
      idata_72_pt_V   : in  std_logic_vector (3 downto 0);
      idata_73_pt_V   : in  std_logic_vector (3 downto 0);
      idata_74_pt_V   : in  std_logic_vector (3 downto 0);
      idata_75_pt_V   : in  std_logic_vector (3 downto 0);
      idata_76_pt_V   : in  std_logic_vector (3 downto 0);
      idata_77_pt_V   : in  std_logic_vector (3 downto 0);
      idata_78_pt_V   : in  std_logic_vector (3 downto 0);
      idata_79_pt_V   : in  std_logic_vector (3 downto 0);
      idata_80_pt_V   : in  std_logic_vector (3 downto 0);
      idata_81_pt_V   : in  std_logic_vector (3 downto 0);
      idata_82_pt_V   : in  std_logic_vector (3 downto 0);
      idata_83_pt_V   : in  std_logic_vector (3 downto 0);
      idata_84_pt_V   : in  std_logic_vector (3 downto 0);
      idata_85_pt_V   : in  std_logic_vector (3 downto 0);
      idata_86_pt_V   : in  std_logic_vector (3 downto 0);
      idata_87_pt_V   : in  std_logic_vector (3 downto 0);
      idata_88_pt_V   : in  std_logic_vector (3 downto 0);
      idata_89_pt_V   : in  std_logic_vector (3 downto 0);
      idata_90_pt_V   : in  std_logic_vector (3 downto 0);
      idata_91_pt_V   : in  std_logic_vector (3 downto 0);
      idata_92_pt_V   : in  std_logic_vector (3 downto 0);
      idata_93_pt_V   : in  std_logic_vector (3 downto 0);
      idata_94_pt_V   : in  std_logic_vector (3 downto 0);
      idata_95_pt_V   : in  std_logic_vector (3 downto 0);
      idata_96_pt_V   : in  std_logic_vector (3 downto 0);
      idata_97_pt_V   : in  std_logic_vector (3 downto 0);
      idata_98_pt_V   : in  std_logic_vector (3 downto 0);
      idata_99_pt_V   : in  std_logic_vector (3 downto 0);
      idata_100_pt_V  : in  std_logic_vector (3 downto 0);
      idata_101_pt_V  : in  std_logic_vector (3 downto 0);
      idata_102_pt_V  : in  std_logic_vector (3 downto 0);
      idata_103_pt_V  : in  std_logic_vector (3 downto 0);
      idata_104_pt_V  : in  std_logic_vector (3 downto 0);
      idata_105_pt_V  : in  std_logic_vector (3 downto 0);
      idata_106_pt_V  : in  std_logic_vector (3 downto 0);
      idata_107_pt_V  : in  std_logic_vector (3 downto 0);
      idata_108_pt_V  : in  std_logic_vector (3 downto 0);
      idata_109_pt_V  : in  std_logic_vector (3 downto 0);
      idata_110_pt_V  : in  std_logic_vector (3 downto 0);
      idata_111_pt_V  : in  std_logic_vector (3 downto 0);
      idata_112_pt_V  : in  std_logic_vector (3 downto 0);
      idata_113_pt_V  : in  std_logic_vector (3 downto 0);
      idata_114_pt_V  : in  std_logic_vector (3 downto 0);
      idata_115_pt_V  : in  std_logic_vector (3 downto 0);
      idata_116_pt_V  : in  std_logic_vector (3 downto 0);
      idata_117_pt_V  : in  std_logic_vector (3 downto 0);
      idata_118_pt_V  : in  std_logic_vector (3 downto 0);
      idata_119_pt_V  : in  std_logic_vector (3 downto 0);
      idata_120_pt_V  : in  std_logic_vector (3 downto 0);
      idata_121_pt_V  : in  std_logic_vector (3 downto 0);
      idata_122_pt_V  : in  std_logic_vector (3 downto 0);
      idata_123_pt_V  : in  std_logic_vector (3 downto 0);
      idata_124_pt_V  : in  std_logic_vector (3 downto 0);
      idata_125_pt_V  : in  std_logic_vector (3 downto 0);
      idata_126_pt_V  : in  std_logic_vector (3 downto 0);
      idata_127_pt_V  : in  std_logic_vector (3 downto 0);
      idata_128_pt_V  : in  std_logic_vector (3 downto 0);
      idata_129_pt_V  : in  std_logic_vector (3 downto 0);
      idata_130_pt_V  : in  std_logic_vector (3 downto 0);
      idata_131_pt_V  : in  std_logic_vector (3 downto 0);
      idata_132_pt_V  : in  std_logic_vector (3 downto 0);
      idata_133_pt_V  : in  std_logic_vector (3 downto 0);
      idata_134_pt_V  : in  std_logic_vector (3 downto 0);
      idata_135_pt_V  : in  std_logic_vector (3 downto 0);
      idata_136_pt_V  : in  std_logic_vector (3 downto 0);
      idata_137_pt_V  : in  std_logic_vector (3 downto 0);
      idata_138_pt_V  : in  std_logic_vector (3 downto 0);
      idata_139_pt_V  : in  std_logic_vector (3 downto 0);
      idata_140_pt_V  : in  std_logic_vector (3 downto 0);
      idata_141_pt_V  : in  std_logic_vector (3 downto 0);
      idata_142_pt_V  : in  std_logic_vector (3 downto 0);
      idata_143_pt_V  : in  std_logic_vector (3 downto 0);
      idata_144_pt_V  : in  std_logic_vector (3 downto 0);
      idata_145_pt_V  : in  std_logic_vector (3 downto 0);
      idata_146_pt_V  : in  std_logic_vector (3 downto 0);
      idata_147_pt_V  : in  std_logic_vector (3 downto 0);
      idata_148_pt_V  : in  std_logic_vector (3 downto 0);
      idata_149_pt_V  : in  std_logic_vector (3 downto 0);
      idata_150_pt_V  : in  std_logic_vector (3 downto 0);
      idata_151_pt_V  : in  std_logic_vector (3 downto 0);
      idata_152_pt_V  : in  std_logic_vector (3 downto 0);
      idata_153_pt_V  : in  std_logic_vector (3 downto 0);
      idata_154_pt_V  : in  std_logic_vector (3 downto 0);
      idata_155_pt_V  : in  std_logic_vector (3 downto 0);
      idata_156_pt_V  : in  std_logic_vector (3 downto 0);
      idata_157_pt_V  : in  std_logic_vector (3 downto 0);
      idata_158_pt_V  : in  std_logic_vector (3 downto 0);
      idata_159_pt_V  : in  std_logic_vector (3 downto 0);
      idata_160_pt_V  : in  std_logic_vector (3 downto 0);
      idata_161_pt_V  : in  std_logic_vector (3 downto 0);
      idata_162_pt_V  : in  std_logic_vector (3 downto 0);
      idata_163_pt_V  : in  std_logic_vector (3 downto 0);
      idata_164_pt_V  : in  std_logic_vector (3 downto 0);
      idata_165_pt_V  : in  std_logic_vector (3 downto 0);
      idata_166_pt_V  : in  std_logic_vector (3 downto 0);
      idata_167_pt_V  : in  std_logic_vector (3 downto 0);
      idata_168_pt_V  : in  std_logic_vector (3 downto 0);
      idata_169_pt_V  : in  std_logic_vector (3 downto 0);
      idata_170_pt_V  : in  std_logic_vector (3 downto 0);
      idata_171_pt_V  : in  std_logic_vector (3 downto 0);
      idata_172_pt_V  : in  std_logic_vector (3 downto 0);
      idata_173_pt_V  : in  std_logic_vector (3 downto 0);
      idata_174_pt_V  : in  std_logic_vector (3 downto 0);
      idata_175_pt_V  : in  std_logic_vector (3 downto 0);
      idata_176_pt_V  : in  std_logic_vector (3 downto 0);
      idata_177_pt_V  : in  std_logic_vector (3 downto 0);
      idata_178_pt_V  : in  std_logic_vector (3 downto 0);
      idata_179_pt_V  : in  std_logic_vector (3 downto 0);
      idata_180_pt_V  : in  std_logic_vector (3 downto 0);
      idata_181_pt_V  : in  std_logic_vector (3 downto 0);
      idata_182_pt_V  : in  std_logic_vector (3 downto 0);
      idata_183_pt_V  : in  std_logic_vector (3 downto 0);
      idata_184_pt_V  : in  std_logic_vector (3 downto 0);
      idata_185_pt_V  : in  std_logic_vector (3 downto 0);
      idata_186_pt_V  : in  std_logic_vector (3 downto 0);
      idata_187_pt_V  : in  std_logic_vector (3 downto 0);
      idata_188_pt_V  : in  std_logic_vector (3 downto 0);
      idata_189_pt_V  : in  std_logic_vector (3 downto 0);
      idata_190_pt_V  : in  std_logic_vector (3 downto 0);
      idata_191_pt_V  : in  std_logic_vector (3 downto 0);
      idata_192_pt_V  : in  std_logic_vector (3 downto 0);
      idata_193_pt_V  : in  std_logic_vector (3 downto 0);
      idata_194_pt_V  : in  std_logic_vector (3 downto 0);
      idata_195_pt_V  : in  std_logic_vector (3 downto 0);
      idata_196_pt_V  : in  std_logic_vector (3 downto 0);
      idata_197_pt_V  : in  std_logic_vector (3 downto 0);
      idata_198_pt_V  : in  std_logic_vector (3 downto 0);
      idata_199_pt_V  : in  std_logic_vector (3 downto 0);
      idata_200_pt_V  : in  std_logic_vector (3 downto 0);
      idata_201_pt_V  : in  std_logic_vector (3 downto 0);
      idata_202_pt_V  : in  std_logic_vector (3 downto 0);
      idata_203_pt_V  : in  std_logic_vector (3 downto 0);
      idata_204_pt_V  : in  std_logic_vector (3 downto 0);
      idata_205_pt_V  : in  std_logic_vector (3 downto 0);
      idata_206_pt_V  : in  std_logic_vector (3 downto 0);
      idata_207_pt_V  : in  std_logic_vector (3 downto 0);
      idata_208_pt_V  : in  std_logic_vector (3 downto 0);
      idata_209_pt_V  : in  std_logic_vector (3 downto 0);
      idata_210_pt_V  : in  std_logic_vector (3 downto 0);
      idata_211_pt_V  : in  std_logic_vector (3 downto 0);
      idata_212_pt_V  : in  std_logic_vector (3 downto 0);
      idata_213_pt_V  : in  std_logic_vector (3 downto 0);
      idata_214_pt_V  : in  std_logic_vector (3 downto 0);
      idata_215_pt_V  : in  std_logic_vector (3 downto 0);
      idata_216_pt_V  : in  std_logic_vector (3 downto 0);
      idata_217_pt_V  : in  std_logic_vector (3 downto 0);
      idata_218_pt_V  : in  std_logic_vector (3 downto 0);
      idata_219_pt_V  : in  std_logic_vector (3 downto 0);
      idata_220_pt_V  : in  std_logic_vector (3 downto 0);
      idata_221_pt_V  : in  std_logic_vector (3 downto 0);
      idata_222_pt_V  : in  std_logic_vector (3 downto 0);
      idata_223_pt_V  : in  std_logic_vector (3 downto 0);
      idata_224_pt_V  : in  std_logic_vector (3 downto 0);
      idata_225_pt_V  : in  std_logic_vector (3 downto 0);
      idata_226_pt_V  : in  std_logic_vector (3 downto 0);
      idata_227_pt_V  : in  std_logic_vector (3 downto 0);
      idata_228_pt_V  : in  std_logic_vector (3 downto 0);
      idata_229_pt_V  : in  std_logic_vector (3 downto 0);
      idata_230_pt_V  : in  std_logic_vector (3 downto 0);
      idata_231_pt_V  : in  std_logic_vector (3 downto 0);
      idata_232_pt_V  : in  std_logic_vector (3 downto 0);
      idata_233_pt_V  : in  std_logic_vector (3 downto 0);
      idata_234_pt_V  : in  std_logic_vector (3 downto 0);
      idata_235_pt_V  : in  std_logic_vector (3 downto 0);
      idata_236_pt_V  : in  std_logic_vector (3 downto 0);
      idata_237_pt_V  : in  std_logic_vector (3 downto 0);
      idata_238_pt_V  : in  std_logic_vector (3 downto 0);
      idata_239_pt_V  : in  std_logic_vector (3 downto 0);
      idata_240_pt_V  : in  std_logic_vector (3 downto 0);
      idata_241_pt_V  : in  std_logic_vector (3 downto 0);
      idata_242_pt_V  : in  std_logic_vector (3 downto 0);
      idata_243_pt_V  : in  std_logic_vector (3 downto 0);
      idata_244_pt_V  : in  std_logic_vector (3 downto 0);
      idata_245_pt_V  : in  std_logic_vector (3 downto 0);
      idata_246_pt_V  : in  std_logic_vector (3 downto 0);
      idata_247_pt_V  : in  std_logic_vector (3 downto 0);
      idata_248_pt_V  : in  std_logic_vector (3 downto 0);
      idata_249_pt_V  : in  std_logic_vector (3 downto 0);
      idata_250_pt_V  : in  std_logic_vector (3 downto 0);
      idata_251_pt_V  : in  std_logic_vector (3 downto 0);
      idata_252_pt_V  : in  std_logic_vector (3 downto 0);
      idata_253_pt_V  : in  std_logic_vector (3 downto 0);
      idata_254_pt_V  : in  std_logic_vector (3 downto 0);
      idata_255_pt_V  : in  std_logic_vector (3 downto 0);
      idata_256_pt_V  : in  std_logic_vector (3 downto 0);
      idata_257_pt_V  : in  std_logic_vector (3 downto 0);
      idata_258_pt_V  : in  std_logic_vector (3 downto 0);
      idata_259_pt_V  : in  std_logic_vector (3 downto 0);
      idata_260_pt_V  : in  std_logic_vector (3 downto 0);
      idata_261_pt_V  : in  std_logic_vector (3 downto 0);
      idata_262_pt_V  : in  std_logic_vector (3 downto 0);
      idata_263_pt_V  : in  std_logic_vector (3 downto 0);
      idata_264_pt_V  : in  std_logic_vector (3 downto 0);
      idata_265_pt_V  : in  std_logic_vector (3 downto 0);
      idata_266_pt_V  : in  std_logic_vector (3 downto 0);
      idata_267_pt_V  : in  std_logic_vector (3 downto 0);
      idata_268_pt_V  : in  std_logic_vector (3 downto 0);
      idata_269_pt_V  : in  std_logic_vector (3 downto 0);
      idata_270_pt_V  : in  std_logic_vector (3 downto 0);
      idata_271_pt_V  : in  std_logic_vector (3 downto 0);
      idata_272_pt_V  : in  std_logic_vector (3 downto 0);
      idata_273_pt_V  : in  std_logic_vector (3 downto 0);
      idata_274_pt_V  : in  std_logic_vector (3 downto 0);
      idata_275_pt_V  : in  std_logic_vector (3 downto 0);
      idata_276_pt_V  : in  std_logic_vector (3 downto 0);
      idata_277_pt_V  : in  std_logic_vector (3 downto 0);
      idata_278_pt_V  : in  std_logic_vector (3 downto 0);
      idata_279_pt_V  : in  std_logic_vector (3 downto 0);
      idata_280_pt_V  : in  std_logic_vector (3 downto 0);
      idata_281_pt_V  : in  std_logic_vector (3 downto 0);
      idata_282_pt_V  : in  std_logic_vector (3 downto 0);
      idata_283_pt_V  : in  std_logic_vector (3 downto 0);
      idata_284_pt_V  : in  std_logic_vector (3 downto 0);
      idata_285_pt_V  : in  std_logic_vector (3 downto 0);
      idata_286_pt_V  : in  std_logic_vector (3 downto 0);
      idata_287_pt_V  : in  std_logic_vector (3 downto 0);
      idata_288_pt_V  : in  std_logic_vector (3 downto 0);
      idata_289_pt_V  : in  std_logic_vector (3 downto 0);
      idata_290_pt_V  : in  std_logic_vector (3 downto 0);
      idata_291_pt_V  : in  std_logic_vector (3 downto 0);
      idata_292_pt_V  : in  std_logic_vector (3 downto 0);
      idata_293_pt_V  : in  std_logic_vector (3 downto 0);
      idata_294_pt_V  : in  std_logic_vector (3 downto 0);
      idata_295_pt_V  : in  std_logic_vector (3 downto 0);
      idata_296_pt_V  : in  std_logic_vector (3 downto 0);
      idata_297_pt_V  : in  std_logic_vector (3 downto 0);
      idata_298_pt_V  : in  std_logic_vector (3 downto 0);
      idata_299_pt_V  : in  std_logic_vector (3 downto 0);
      idata_300_pt_V  : in  std_logic_vector (3 downto 0);
      idata_301_pt_V  : in  std_logic_vector (3 downto 0);
      idata_302_pt_V  : in  std_logic_vector (3 downto 0);
      idata_303_pt_V  : in  std_logic_vector (3 downto 0);
      idata_304_pt_V  : in  std_logic_vector (3 downto 0);
      idata_305_pt_V  : in  std_logic_vector (3 downto 0);
      idata_306_pt_V  : in  std_logic_vector (3 downto 0);
      idata_307_pt_V  : in  std_logic_vector (3 downto 0);
      idata_308_pt_V  : in  std_logic_vector (3 downto 0);
      idata_309_pt_V  : in  std_logic_vector (3 downto 0);
      idata_310_pt_V  : in  std_logic_vector (3 downto 0);
      idata_311_pt_V  : in  std_logic_vector (3 downto 0);
      idata_312_pt_V  : in  std_logic_vector (3 downto 0);
      idata_313_pt_V  : in  std_logic_vector (3 downto 0);
      idata_314_pt_V  : in  std_logic_vector (3 downto 0);
      idata_315_pt_V  : in  std_logic_vector (3 downto 0);
      idata_316_pt_V  : in  std_logic_vector (3 downto 0);
      idata_317_pt_V  : in  std_logic_vector (3 downto 0);
      idata_318_pt_V  : in  std_logic_vector (3 downto 0);
      idata_319_pt_V  : in  std_logic_vector (3 downto 0);
      idata_320_pt_V  : in  std_logic_vector (3 downto 0);
      idata_321_pt_V  : in  std_logic_vector (3 downto 0);
      idata_322_pt_V  : in  std_logic_vector (3 downto 0);
      idata_323_pt_V  : in  std_logic_vector (3 downto 0);
      idata_324_pt_V  : in  std_logic_vector (3 downto 0);
      idata_325_pt_V  : in  std_logic_vector (3 downto 0);
      idata_326_pt_V  : in  std_logic_vector (3 downto 0);
      idata_327_pt_V  : in  std_logic_vector (3 downto 0);
      idata_328_pt_V  : in  std_logic_vector (3 downto 0);
      idata_329_pt_V  : in  std_logic_vector (3 downto 0);
      idata_330_pt_V  : in  std_logic_vector (3 downto 0);
      idata_331_pt_V  : in  std_logic_vector (3 downto 0);
      idata_332_pt_V  : in  std_logic_vector (3 downto 0);
      idata_333_pt_V  : in  std_logic_vector (3 downto 0);
      idata_334_pt_V  : in  std_logic_vector (3 downto 0);
      idata_335_pt_V  : in  std_logic_vector (3 downto 0);
      idata_336_pt_V  : in  std_logic_vector (3 downto 0);
      idata_337_pt_V  : in  std_logic_vector (3 downto 0);
      idata_338_pt_V  : in  std_logic_vector (3 downto 0);
      idata_339_pt_V  : in  std_logic_vector (3 downto 0);
      idata_340_pt_V  : in  std_logic_vector (3 downto 0);
      idata_341_pt_V  : in  std_logic_vector (3 downto 0);
      idata_342_pt_V  : in  std_logic_vector (3 downto 0);
      idata_343_pt_V  : in  std_logic_vector (3 downto 0);
      idata_344_pt_V  : in  std_logic_vector (3 downto 0);
      idata_345_pt_V  : in  std_logic_vector (3 downto 0);
      idata_346_pt_V  : in  std_logic_vector (3 downto 0);
      idata_347_pt_V  : in  std_logic_vector (3 downto 0);
      idata_348_pt_V  : in  std_logic_vector (3 downto 0);
      idata_349_pt_V  : in  std_logic_vector (3 downto 0);
      idata_350_pt_V  : in  std_logic_vector (3 downto 0);
      idata_351_pt_V  : in  std_logic_vector (3 downto 0);
      idata_0_roi_V   : in  std_logic_vector (7 downto 0);
      idata_1_roi_V   : in  std_logic_vector (7 downto 0);
      idata_2_roi_V   : in  std_logic_vector (7 downto 0);
      idata_3_roi_V   : in  std_logic_vector (7 downto 0);
      idata_4_roi_V   : in  std_logic_vector (7 downto 0);
      idata_5_roi_V   : in  std_logic_vector (7 downto 0);
      idata_6_roi_V   : in  std_logic_vector (7 downto 0);
      idata_7_roi_V   : in  std_logic_vector (7 downto 0);
      idata_8_roi_V   : in  std_logic_vector (7 downto 0);
      idata_9_roi_V   : in  std_logic_vector (7 downto 0);
      idata_10_roi_V  : in  std_logic_vector (7 downto 0);
      idata_11_roi_V  : in  std_logic_vector (7 downto 0);
      idata_12_roi_V  : in  std_logic_vector (7 downto 0);
      idata_13_roi_V  : in  std_logic_vector (7 downto 0);
      idata_14_roi_V  : in  std_logic_vector (7 downto 0);
      idata_15_roi_V  : in  std_logic_vector (7 downto 0);
      idata_16_roi_V  : in  std_logic_vector (7 downto 0);
      idata_17_roi_V  : in  std_logic_vector (7 downto 0);
      idata_18_roi_V  : in  std_logic_vector (7 downto 0);
      idata_19_roi_V  : in  std_logic_vector (7 downto 0);
      idata_20_roi_V  : in  std_logic_vector (7 downto 0);
      idata_21_roi_V  : in  std_logic_vector (7 downto 0);
      idata_22_roi_V  : in  std_logic_vector (7 downto 0);
      idata_23_roi_V  : in  std_logic_vector (7 downto 0);
      idata_24_roi_V  : in  std_logic_vector (7 downto 0);
      idata_25_roi_V  : in  std_logic_vector (7 downto 0);
      idata_26_roi_V  : in  std_logic_vector (7 downto 0);
      idata_27_roi_V  : in  std_logic_vector (7 downto 0);
      idata_28_roi_V  : in  std_logic_vector (7 downto 0);
      idata_29_roi_V  : in  std_logic_vector (7 downto 0);
      idata_30_roi_V  : in  std_logic_vector (7 downto 0);
      idata_31_roi_V  : in  std_logic_vector (7 downto 0);
      idata_32_roi_V  : in  std_logic_vector (7 downto 0);
      idata_33_roi_V  : in  std_logic_vector (7 downto 0);
      idata_34_roi_V  : in  std_logic_vector (7 downto 0);
      idata_35_roi_V  : in  std_logic_vector (7 downto 0);
      idata_36_roi_V  : in  std_logic_vector (7 downto 0);
      idata_37_roi_V  : in  std_logic_vector (7 downto 0);
      idata_38_roi_V  : in  std_logic_vector (7 downto 0);
      idata_39_roi_V  : in  std_logic_vector (7 downto 0);
      idata_40_roi_V  : in  std_logic_vector (7 downto 0);
      idata_41_roi_V  : in  std_logic_vector (7 downto 0);
      idata_42_roi_V  : in  std_logic_vector (7 downto 0);
      idata_43_roi_V  : in  std_logic_vector (7 downto 0);
      idata_44_roi_V  : in  std_logic_vector (7 downto 0);
      idata_45_roi_V  : in  std_logic_vector (7 downto 0);
      idata_46_roi_V  : in  std_logic_vector (7 downto 0);
      idata_47_roi_V  : in  std_logic_vector (7 downto 0);
      idata_48_roi_V  : in  std_logic_vector (7 downto 0);
      idata_49_roi_V  : in  std_logic_vector (7 downto 0);
      idata_50_roi_V  : in  std_logic_vector (7 downto 0);
      idata_51_roi_V  : in  std_logic_vector (7 downto 0);
      idata_52_roi_V  : in  std_logic_vector (7 downto 0);
      idata_53_roi_V  : in  std_logic_vector (7 downto 0);
      idata_54_roi_V  : in  std_logic_vector (7 downto 0);
      idata_55_roi_V  : in  std_logic_vector (7 downto 0);
      idata_56_roi_V  : in  std_logic_vector (7 downto 0);
      idata_57_roi_V  : in  std_logic_vector (7 downto 0);
      idata_58_roi_V  : in  std_logic_vector (7 downto 0);
      idata_59_roi_V  : in  std_logic_vector (7 downto 0);
      idata_60_roi_V  : in  std_logic_vector (7 downto 0);
      idata_61_roi_V  : in  std_logic_vector (7 downto 0);
      idata_62_roi_V  : in  std_logic_vector (7 downto 0);
      idata_63_roi_V  : in  std_logic_vector (7 downto 0);
      idata_64_roi_V  : in  std_logic_vector (7 downto 0);
      idata_65_roi_V  : in  std_logic_vector (7 downto 0);
      idata_66_roi_V  : in  std_logic_vector (7 downto 0);
      idata_67_roi_V  : in  std_logic_vector (7 downto 0);
      idata_68_roi_V  : in  std_logic_vector (7 downto 0);
      idata_69_roi_V  : in  std_logic_vector (7 downto 0);
      idata_70_roi_V  : in  std_logic_vector (7 downto 0);
      idata_71_roi_V  : in  std_logic_vector (7 downto 0);
      idata_72_roi_V  : in  std_logic_vector (7 downto 0);
      idata_73_roi_V  : in  std_logic_vector (7 downto 0);
      idata_74_roi_V  : in  std_logic_vector (7 downto 0);
      idata_75_roi_V  : in  std_logic_vector (7 downto 0);
      idata_76_roi_V  : in  std_logic_vector (7 downto 0);
      idata_77_roi_V  : in  std_logic_vector (7 downto 0);
      idata_78_roi_V  : in  std_logic_vector (7 downto 0);
      idata_79_roi_V  : in  std_logic_vector (7 downto 0);
      idata_80_roi_V  : in  std_logic_vector (7 downto 0);
      idata_81_roi_V  : in  std_logic_vector (7 downto 0);
      idata_82_roi_V  : in  std_logic_vector (7 downto 0);
      idata_83_roi_V  : in  std_logic_vector (7 downto 0);
      idata_84_roi_V  : in  std_logic_vector (7 downto 0);
      idata_85_roi_V  : in  std_logic_vector (7 downto 0);
      idata_86_roi_V  : in  std_logic_vector (7 downto 0);
      idata_87_roi_V  : in  std_logic_vector (7 downto 0);
      idata_88_roi_V  : in  std_logic_vector (7 downto 0);
      idata_89_roi_V  : in  std_logic_vector (7 downto 0);
      idata_90_roi_V  : in  std_logic_vector (7 downto 0);
      idata_91_roi_V  : in  std_logic_vector (7 downto 0);
      idata_92_roi_V  : in  std_logic_vector (7 downto 0);
      idata_93_roi_V  : in  std_logic_vector (7 downto 0);
      idata_94_roi_V  : in  std_logic_vector (7 downto 0);
      idata_95_roi_V  : in  std_logic_vector (7 downto 0);
      idata_96_roi_V  : in  std_logic_vector (7 downto 0);
      idata_97_roi_V  : in  std_logic_vector (7 downto 0);
      idata_98_roi_V  : in  std_logic_vector (7 downto 0);
      idata_99_roi_V  : in  std_logic_vector (7 downto 0);
      idata_100_roi_V : in  std_logic_vector (7 downto 0);
      idata_101_roi_V : in  std_logic_vector (7 downto 0);
      idata_102_roi_V : in  std_logic_vector (7 downto 0);
      idata_103_roi_V : in  std_logic_vector (7 downto 0);
      idata_104_roi_V : in  std_logic_vector (7 downto 0);
      idata_105_roi_V : in  std_logic_vector (7 downto 0);
      idata_106_roi_V : in  std_logic_vector (7 downto 0);
      idata_107_roi_V : in  std_logic_vector (7 downto 0);
      idata_108_roi_V : in  std_logic_vector (7 downto 0);
      idata_109_roi_V : in  std_logic_vector (7 downto 0);
      idata_110_roi_V : in  std_logic_vector (7 downto 0);
      idata_111_roi_V : in  std_logic_vector (7 downto 0);
      idata_112_roi_V : in  std_logic_vector (7 downto 0);
      idata_113_roi_V : in  std_logic_vector (7 downto 0);
      idata_114_roi_V : in  std_logic_vector (7 downto 0);
      idata_115_roi_V : in  std_logic_vector (7 downto 0);
      idata_116_roi_V : in  std_logic_vector (7 downto 0);
      idata_117_roi_V : in  std_logic_vector (7 downto 0);
      idata_118_roi_V : in  std_logic_vector (7 downto 0);
      idata_119_roi_V : in  std_logic_vector (7 downto 0);
      idata_120_roi_V : in  std_logic_vector (7 downto 0);
      idata_121_roi_V : in  std_logic_vector (7 downto 0);
      idata_122_roi_V : in  std_logic_vector (7 downto 0);
      idata_123_roi_V : in  std_logic_vector (7 downto 0);
      idata_124_roi_V : in  std_logic_vector (7 downto 0);
      idata_125_roi_V : in  std_logic_vector (7 downto 0);
      idata_126_roi_V : in  std_logic_vector (7 downto 0);
      idata_127_roi_V : in  std_logic_vector (7 downto 0);
      idata_128_roi_V : in  std_logic_vector (7 downto 0);
      idata_129_roi_V : in  std_logic_vector (7 downto 0);
      idata_130_roi_V : in  std_logic_vector (7 downto 0);
      idata_131_roi_V : in  std_logic_vector (7 downto 0);
      idata_132_roi_V : in  std_logic_vector (7 downto 0);
      idata_133_roi_V : in  std_logic_vector (7 downto 0);
      idata_134_roi_V : in  std_logic_vector (7 downto 0);
      idata_135_roi_V : in  std_logic_vector (7 downto 0);
      idata_136_roi_V : in  std_logic_vector (7 downto 0);
      idata_137_roi_V : in  std_logic_vector (7 downto 0);
      idata_138_roi_V : in  std_logic_vector (7 downto 0);
      idata_139_roi_V : in  std_logic_vector (7 downto 0);
      idata_140_roi_V : in  std_logic_vector (7 downto 0);
      idata_141_roi_V : in  std_logic_vector (7 downto 0);
      idata_142_roi_V : in  std_logic_vector (7 downto 0);
      idata_143_roi_V : in  std_logic_vector (7 downto 0);
      idata_144_roi_V : in  std_logic_vector (7 downto 0);
      idata_145_roi_V : in  std_logic_vector (7 downto 0);
      idata_146_roi_V : in  std_logic_vector (7 downto 0);
      idata_147_roi_V : in  std_logic_vector (7 downto 0);
      idata_148_roi_V : in  std_logic_vector (7 downto 0);
      idata_149_roi_V : in  std_logic_vector (7 downto 0);
      idata_150_roi_V : in  std_logic_vector (7 downto 0);
      idata_151_roi_V : in  std_logic_vector (7 downto 0);
      idata_152_roi_V : in  std_logic_vector (7 downto 0);
      idata_153_roi_V : in  std_logic_vector (7 downto 0);
      idata_154_roi_V : in  std_logic_vector (7 downto 0);
      idata_155_roi_V : in  std_logic_vector (7 downto 0);
      idata_156_roi_V : in  std_logic_vector (7 downto 0);
      idata_157_roi_V : in  std_logic_vector (7 downto 0);
      idata_158_roi_V : in  std_logic_vector (7 downto 0);
      idata_159_roi_V : in  std_logic_vector (7 downto 0);
      idata_160_roi_V : in  std_logic_vector (7 downto 0);
      idata_161_roi_V : in  std_logic_vector (7 downto 0);
      idata_162_roi_V : in  std_logic_vector (7 downto 0);
      idata_163_roi_V : in  std_logic_vector (7 downto 0);
      idata_164_roi_V : in  std_logic_vector (7 downto 0);
      idata_165_roi_V : in  std_logic_vector (7 downto 0);
      idata_166_roi_V : in  std_logic_vector (7 downto 0);
      idata_167_roi_V : in  std_logic_vector (7 downto 0);
      idata_168_roi_V : in  std_logic_vector (7 downto 0);
      idata_169_roi_V : in  std_logic_vector (7 downto 0);
      idata_170_roi_V : in  std_logic_vector (7 downto 0);
      idata_171_roi_V : in  std_logic_vector (7 downto 0);
      idata_172_roi_V : in  std_logic_vector (7 downto 0);
      idata_173_roi_V : in  std_logic_vector (7 downto 0);
      idata_174_roi_V : in  std_logic_vector (7 downto 0);
      idata_175_roi_V : in  std_logic_vector (7 downto 0);
      idata_176_roi_V : in  std_logic_vector (7 downto 0);
      idata_177_roi_V : in  std_logic_vector (7 downto 0);
      idata_178_roi_V : in  std_logic_vector (7 downto 0);
      idata_179_roi_V : in  std_logic_vector (7 downto 0);
      idata_180_roi_V : in  std_logic_vector (7 downto 0);
      idata_181_roi_V : in  std_logic_vector (7 downto 0);
      idata_182_roi_V : in  std_logic_vector (7 downto 0);
      idata_183_roi_V : in  std_logic_vector (7 downto 0);
      idata_184_roi_V : in  std_logic_vector (7 downto 0);
      idata_185_roi_V : in  std_logic_vector (7 downto 0);
      idata_186_roi_V : in  std_logic_vector (7 downto 0);
      idata_187_roi_V : in  std_logic_vector (7 downto 0);
      idata_188_roi_V : in  std_logic_vector (7 downto 0);
      idata_189_roi_V : in  std_logic_vector (7 downto 0);
      idata_190_roi_V : in  std_logic_vector (7 downto 0);
      idata_191_roi_V : in  std_logic_vector (7 downto 0);
      idata_192_roi_V : in  std_logic_vector (7 downto 0);
      idata_193_roi_V : in  std_logic_vector (7 downto 0);
      idata_194_roi_V : in  std_logic_vector (7 downto 0);
      idata_195_roi_V : in  std_logic_vector (7 downto 0);
      idata_196_roi_V : in  std_logic_vector (7 downto 0);
      idata_197_roi_V : in  std_logic_vector (7 downto 0);
      idata_198_roi_V : in  std_logic_vector (7 downto 0);
      idata_199_roi_V : in  std_logic_vector (7 downto 0);
      idata_200_roi_V : in  std_logic_vector (7 downto 0);
      idata_201_roi_V : in  std_logic_vector (7 downto 0);
      idata_202_roi_V : in  std_logic_vector (7 downto 0);
      idata_203_roi_V : in  std_logic_vector (7 downto 0);
      idata_204_roi_V : in  std_logic_vector (7 downto 0);
      idata_205_roi_V : in  std_logic_vector (7 downto 0);
      idata_206_roi_V : in  std_logic_vector (7 downto 0);
      idata_207_roi_V : in  std_logic_vector (7 downto 0);
      idata_208_roi_V : in  std_logic_vector (7 downto 0);
      idata_209_roi_V : in  std_logic_vector (7 downto 0);
      idata_210_roi_V : in  std_logic_vector (7 downto 0);
      idata_211_roi_V : in  std_logic_vector (7 downto 0);
      idata_212_roi_V : in  std_logic_vector (7 downto 0);
      idata_213_roi_V : in  std_logic_vector (7 downto 0);
      idata_214_roi_V : in  std_logic_vector (7 downto 0);
      idata_215_roi_V : in  std_logic_vector (7 downto 0);
      idata_216_roi_V : in  std_logic_vector (7 downto 0);
      idata_217_roi_V : in  std_logic_vector (7 downto 0);
      idata_218_roi_V : in  std_logic_vector (7 downto 0);
      idata_219_roi_V : in  std_logic_vector (7 downto 0);
      idata_220_roi_V : in  std_logic_vector (7 downto 0);
      idata_221_roi_V : in  std_logic_vector (7 downto 0);
      idata_222_roi_V : in  std_logic_vector (7 downto 0);
      idata_223_roi_V : in  std_logic_vector (7 downto 0);
      idata_224_roi_V : in  std_logic_vector (7 downto 0);
      idata_225_roi_V : in  std_logic_vector (7 downto 0);
      idata_226_roi_V : in  std_logic_vector (7 downto 0);
      idata_227_roi_V : in  std_logic_vector (7 downto 0);
      idata_228_roi_V : in  std_logic_vector (7 downto 0);
      idata_229_roi_V : in  std_logic_vector (7 downto 0);
      idata_230_roi_V : in  std_logic_vector (7 downto 0);
      idata_231_roi_V : in  std_logic_vector (7 downto 0);
      idata_232_roi_V : in  std_logic_vector (7 downto 0);
      idata_233_roi_V : in  std_logic_vector (7 downto 0);
      idata_234_roi_V : in  std_logic_vector (7 downto 0);
      idata_235_roi_V : in  std_logic_vector (7 downto 0);
      idata_236_roi_V : in  std_logic_vector (7 downto 0);
      idata_237_roi_V : in  std_logic_vector (7 downto 0);
      idata_238_roi_V : in  std_logic_vector (7 downto 0);
      idata_239_roi_V : in  std_logic_vector (7 downto 0);
      idata_240_roi_V : in  std_logic_vector (7 downto 0);
      idata_241_roi_V : in  std_logic_vector (7 downto 0);
      idata_242_roi_V : in  std_logic_vector (7 downto 0);
      idata_243_roi_V : in  std_logic_vector (7 downto 0);
      idata_244_roi_V : in  std_logic_vector (7 downto 0);
      idata_245_roi_V : in  std_logic_vector (7 downto 0);
      idata_246_roi_V : in  std_logic_vector (7 downto 0);
      idata_247_roi_V : in  std_logic_vector (7 downto 0);
      idata_248_roi_V : in  std_logic_vector (7 downto 0);
      idata_249_roi_V : in  std_logic_vector (7 downto 0);
      idata_250_roi_V : in  std_logic_vector (7 downto 0);
      idata_251_roi_V : in  std_logic_vector (7 downto 0);
      idata_252_roi_V : in  std_logic_vector (7 downto 0);
      idata_253_roi_V : in  std_logic_vector (7 downto 0);
      idata_254_roi_V : in  std_logic_vector (7 downto 0);
      idata_255_roi_V : in  std_logic_vector (7 downto 0);
      idata_256_roi_V : in  std_logic_vector (7 downto 0);
      idata_257_roi_V : in  std_logic_vector (7 downto 0);
      idata_258_roi_V : in  std_logic_vector (7 downto 0);
      idata_259_roi_V : in  std_logic_vector (7 downto 0);
      idata_260_roi_V : in  std_logic_vector (7 downto 0);
      idata_261_roi_V : in  std_logic_vector (7 downto 0);
      idata_262_roi_V : in  std_logic_vector (7 downto 0);
      idata_263_roi_V : in  std_logic_vector (7 downto 0);
      idata_264_roi_V : in  std_logic_vector (7 downto 0);
      idata_265_roi_V : in  std_logic_vector (7 downto 0);
      idata_266_roi_V : in  std_logic_vector (7 downto 0);
      idata_267_roi_V : in  std_logic_vector (7 downto 0);
      idata_268_roi_V : in  std_logic_vector (7 downto 0);
      idata_269_roi_V : in  std_logic_vector (7 downto 0);
      idata_270_roi_V : in  std_logic_vector (7 downto 0);
      idata_271_roi_V : in  std_logic_vector (7 downto 0);
      idata_272_roi_V : in  std_logic_vector (7 downto 0);
      idata_273_roi_V : in  std_logic_vector (7 downto 0);
      idata_274_roi_V : in  std_logic_vector (7 downto 0);
      idata_275_roi_V : in  std_logic_vector (7 downto 0);
      idata_276_roi_V : in  std_logic_vector (7 downto 0);
      idata_277_roi_V : in  std_logic_vector (7 downto 0);
      idata_278_roi_V : in  std_logic_vector (7 downto 0);
      idata_279_roi_V : in  std_logic_vector (7 downto 0);
      idata_280_roi_V : in  std_logic_vector (7 downto 0);
      idata_281_roi_V : in  std_logic_vector (7 downto 0);
      idata_282_roi_V : in  std_logic_vector (7 downto 0);
      idata_283_roi_V : in  std_logic_vector (7 downto 0);
      idata_284_roi_V : in  std_logic_vector (7 downto 0);
      idata_285_roi_V : in  std_logic_vector (7 downto 0);
      idata_286_roi_V : in  std_logic_vector (7 downto 0);
      idata_287_roi_V : in  std_logic_vector (7 downto 0);
      idata_288_roi_V : in  std_logic_vector (7 downto 0);
      idata_289_roi_V : in  std_logic_vector (7 downto 0);
      idata_290_roi_V : in  std_logic_vector (7 downto 0);
      idata_291_roi_V : in  std_logic_vector (7 downto 0);
      idata_292_roi_V : in  std_logic_vector (7 downto 0);
      idata_293_roi_V : in  std_logic_vector (7 downto 0);
      idata_294_roi_V : in  std_logic_vector (7 downto 0);
      idata_295_roi_V : in  std_logic_vector (7 downto 0);
      idata_296_roi_V : in  std_logic_vector (7 downto 0);
      idata_297_roi_V : in  std_logic_vector (7 downto 0);
      idata_298_roi_V : in  std_logic_vector (7 downto 0);
      idata_299_roi_V : in  std_logic_vector (7 downto 0);
      idata_300_roi_V : in  std_logic_vector (7 downto 0);
      idata_301_roi_V : in  std_logic_vector (7 downto 0);
      idata_302_roi_V : in  std_logic_vector (7 downto 0);
      idata_303_roi_V : in  std_logic_vector (7 downto 0);
      idata_304_roi_V : in  std_logic_vector (7 downto 0);
      idata_305_roi_V : in  std_logic_vector (7 downto 0);
      idata_306_roi_V : in  std_logic_vector (7 downto 0);
      idata_307_roi_V : in  std_logic_vector (7 downto 0);
      idata_308_roi_V : in  std_logic_vector (7 downto 0);
      idata_309_roi_V : in  std_logic_vector (7 downto 0);
      idata_310_roi_V : in  std_logic_vector (7 downto 0);
      idata_311_roi_V : in  std_logic_vector (7 downto 0);
      idata_312_roi_V : in  std_logic_vector (7 downto 0);
      idata_313_roi_V : in  std_logic_vector (7 downto 0);
      idata_314_roi_V : in  std_logic_vector (7 downto 0);
      idata_315_roi_V : in  std_logic_vector (7 downto 0);
      idata_316_roi_V : in  std_logic_vector (7 downto 0);
      idata_317_roi_V : in  std_logic_vector (7 downto 0);
      idata_318_roi_V : in  std_logic_vector (7 downto 0);
      idata_319_roi_V : in  std_logic_vector (7 downto 0);
      idata_320_roi_V : in  std_logic_vector (7 downto 0);
      idata_321_roi_V : in  std_logic_vector (7 downto 0);
      idata_322_roi_V : in  std_logic_vector (7 downto 0);
      idata_323_roi_V : in  std_logic_vector (7 downto 0);
      idata_324_roi_V : in  std_logic_vector (7 downto 0);
      idata_325_roi_V : in  std_logic_vector (7 downto 0);
      idata_326_roi_V : in  std_logic_vector (7 downto 0);
      idata_327_roi_V : in  std_logic_vector (7 downto 0);
      idata_328_roi_V : in  std_logic_vector (7 downto 0);
      idata_329_roi_V : in  std_logic_vector (7 downto 0);
      idata_330_roi_V : in  std_logic_vector (7 downto 0);
      idata_331_roi_V : in  std_logic_vector (7 downto 0);
      idata_332_roi_V : in  std_logic_vector (7 downto 0);
      idata_333_roi_V : in  std_logic_vector (7 downto 0);
      idata_334_roi_V : in  std_logic_vector (7 downto 0);
      idata_335_roi_V : in  std_logic_vector (7 downto 0);
      idata_336_roi_V : in  std_logic_vector (7 downto 0);
      idata_337_roi_V : in  std_logic_vector (7 downto 0);
      idata_338_roi_V : in  std_logic_vector (7 downto 0);
      idata_339_roi_V : in  std_logic_vector (7 downto 0);
      idata_340_roi_V : in  std_logic_vector (7 downto 0);
      idata_341_roi_V : in  std_logic_vector (7 downto 0);
      idata_342_roi_V : in  std_logic_vector (7 downto 0);
      idata_343_roi_V : in  std_logic_vector (7 downto 0);
      idata_344_roi_V : in  std_logic_vector (7 downto 0);
      idata_345_roi_V : in  std_logic_vector (7 downto 0);
      idata_346_roi_V : in  std_logic_vector (7 downto 0);
      idata_347_roi_V : in  std_logic_vector (7 downto 0);
      idata_348_roi_V : in  std_logic_vector (7 downto 0);
      idata_349_roi_V : in  std_logic_vector (7 downto 0);
      idata_350_roi_V : in  std_logic_vector (7 downto 0);
      idata_351_roi_V : in  std_logic_vector (7 downto 0);
      idata_0_flg_V   : in  std_logic_vector (3 downto 0);
      idata_1_flg_V   : in  std_logic_vector (3 downto 0);
      idata_2_flg_V   : in  std_logic_vector (3 downto 0);
      idata_3_flg_V   : in  std_logic_vector (3 downto 0);
      idata_4_flg_V   : in  std_logic_vector (3 downto 0);
      idata_5_flg_V   : in  std_logic_vector (3 downto 0);
      idata_6_flg_V   : in  std_logic_vector (3 downto 0);
      idata_7_flg_V   : in  std_logic_vector (3 downto 0);
      idata_8_flg_V   : in  std_logic_vector (3 downto 0);
      idata_9_flg_V   : in  std_logic_vector (3 downto 0);
      idata_10_flg_V  : in  std_logic_vector (3 downto 0);
      idata_11_flg_V  : in  std_logic_vector (3 downto 0);
      idata_12_flg_V  : in  std_logic_vector (3 downto 0);
      idata_13_flg_V  : in  std_logic_vector (3 downto 0);
      idata_14_flg_V  : in  std_logic_vector (3 downto 0);
      idata_15_flg_V  : in  std_logic_vector (3 downto 0);
      idata_16_flg_V  : in  std_logic_vector (3 downto 0);
      idata_17_flg_V  : in  std_logic_vector (3 downto 0);
      idata_18_flg_V  : in  std_logic_vector (3 downto 0);
      idata_19_flg_V  : in  std_logic_vector (3 downto 0);
      idata_20_flg_V  : in  std_logic_vector (3 downto 0);
      idata_21_flg_V  : in  std_logic_vector (3 downto 0);
      idata_22_flg_V  : in  std_logic_vector (3 downto 0);
      idata_23_flg_V  : in  std_logic_vector (3 downto 0);
      idata_24_flg_V  : in  std_logic_vector (3 downto 0);
      idata_25_flg_V  : in  std_logic_vector (3 downto 0);
      idata_26_flg_V  : in  std_logic_vector (3 downto 0);
      idata_27_flg_V  : in  std_logic_vector (3 downto 0);
      idata_28_flg_V  : in  std_logic_vector (3 downto 0);
      idata_29_flg_V  : in  std_logic_vector (3 downto 0);
      idata_30_flg_V  : in  std_logic_vector (3 downto 0);
      idata_31_flg_V  : in  std_logic_vector (3 downto 0);
      idata_32_flg_V  : in  std_logic_vector (3 downto 0);
      idata_33_flg_V  : in  std_logic_vector (3 downto 0);
      idata_34_flg_V  : in  std_logic_vector (3 downto 0);
      idata_35_flg_V  : in  std_logic_vector (3 downto 0);
      idata_36_flg_V  : in  std_logic_vector (3 downto 0);
      idata_37_flg_V  : in  std_logic_vector (3 downto 0);
      idata_38_flg_V  : in  std_logic_vector (3 downto 0);
      idata_39_flg_V  : in  std_logic_vector (3 downto 0);
      idata_40_flg_V  : in  std_logic_vector (3 downto 0);
      idata_41_flg_V  : in  std_logic_vector (3 downto 0);
      idata_42_flg_V  : in  std_logic_vector (3 downto 0);
      idata_43_flg_V  : in  std_logic_vector (3 downto 0);
      idata_44_flg_V  : in  std_logic_vector (3 downto 0);
      idata_45_flg_V  : in  std_logic_vector (3 downto 0);
      idata_46_flg_V  : in  std_logic_vector (3 downto 0);
      idata_47_flg_V  : in  std_logic_vector (3 downto 0);
      idata_48_flg_V  : in  std_logic_vector (3 downto 0);
      idata_49_flg_V  : in  std_logic_vector (3 downto 0);
      idata_50_flg_V  : in  std_logic_vector (3 downto 0);
      idata_51_flg_V  : in  std_logic_vector (3 downto 0);
      idata_52_flg_V  : in  std_logic_vector (3 downto 0);
      idata_53_flg_V  : in  std_logic_vector (3 downto 0);
      idata_54_flg_V  : in  std_logic_vector (3 downto 0);
      idata_55_flg_V  : in  std_logic_vector (3 downto 0);
      idata_56_flg_V  : in  std_logic_vector (3 downto 0);
      idata_57_flg_V  : in  std_logic_vector (3 downto 0);
      idata_58_flg_V  : in  std_logic_vector (3 downto 0);
      idata_59_flg_V  : in  std_logic_vector (3 downto 0);
      idata_60_flg_V  : in  std_logic_vector (3 downto 0);
      idata_61_flg_V  : in  std_logic_vector (3 downto 0);
      idata_62_flg_V  : in  std_logic_vector (3 downto 0);
      idata_63_flg_V  : in  std_logic_vector (3 downto 0);
      idata_64_flg_V  : in  std_logic_vector (3 downto 0);
      idata_65_flg_V  : in  std_logic_vector (3 downto 0);
      idata_66_flg_V  : in  std_logic_vector (3 downto 0);
      idata_67_flg_V  : in  std_logic_vector (3 downto 0);
      idata_68_flg_V  : in  std_logic_vector (3 downto 0);
      idata_69_flg_V  : in  std_logic_vector (3 downto 0);
      idata_70_flg_V  : in  std_logic_vector (3 downto 0);
      idata_71_flg_V  : in  std_logic_vector (3 downto 0);
      idata_72_flg_V  : in  std_logic_vector (3 downto 0);
      idata_73_flg_V  : in  std_logic_vector (3 downto 0);
      idata_74_flg_V  : in  std_logic_vector (3 downto 0);
      idata_75_flg_V  : in  std_logic_vector (3 downto 0);
      idata_76_flg_V  : in  std_logic_vector (3 downto 0);
      idata_77_flg_V  : in  std_logic_vector (3 downto 0);
      idata_78_flg_V  : in  std_logic_vector (3 downto 0);
      idata_79_flg_V  : in  std_logic_vector (3 downto 0);
      idata_80_flg_V  : in  std_logic_vector (3 downto 0);
      idata_81_flg_V  : in  std_logic_vector (3 downto 0);
      idata_82_flg_V  : in  std_logic_vector (3 downto 0);
      idata_83_flg_V  : in  std_logic_vector (3 downto 0);
      idata_84_flg_V  : in  std_logic_vector (3 downto 0);
      idata_85_flg_V  : in  std_logic_vector (3 downto 0);
      idata_86_flg_V  : in  std_logic_vector (3 downto 0);
      idata_87_flg_V  : in  std_logic_vector (3 downto 0);
      idata_88_flg_V  : in  std_logic_vector (3 downto 0);
      idata_89_flg_V  : in  std_logic_vector (3 downto 0);
      idata_90_flg_V  : in  std_logic_vector (3 downto 0);
      idata_91_flg_V  : in  std_logic_vector (3 downto 0);
      idata_92_flg_V  : in  std_logic_vector (3 downto 0);
      idata_93_flg_V  : in  std_logic_vector (3 downto 0);
      idata_94_flg_V  : in  std_logic_vector (3 downto 0);
      idata_95_flg_V  : in  std_logic_vector (3 downto 0);
      idata_96_flg_V  : in  std_logic_vector (3 downto 0);
      idata_97_flg_V  : in  std_logic_vector (3 downto 0);
      idata_98_flg_V  : in  std_logic_vector (3 downto 0);
      idata_99_flg_V  : in  std_logic_vector (3 downto 0);
      idata_100_flg_V : in  std_logic_vector (3 downto 0);
      idata_101_flg_V : in  std_logic_vector (3 downto 0);
      idata_102_flg_V : in  std_logic_vector (3 downto 0);
      idata_103_flg_V : in  std_logic_vector (3 downto 0);
      idata_104_flg_V : in  std_logic_vector (3 downto 0);
      idata_105_flg_V : in  std_logic_vector (3 downto 0);
      idata_106_flg_V : in  std_logic_vector (3 downto 0);
      idata_107_flg_V : in  std_logic_vector (3 downto 0);
      idata_108_flg_V : in  std_logic_vector (3 downto 0);
      idata_109_flg_V : in  std_logic_vector (3 downto 0);
      idata_110_flg_V : in  std_logic_vector (3 downto 0);
      idata_111_flg_V : in  std_logic_vector (3 downto 0);
      idata_112_flg_V : in  std_logic_vector (3 downto 0);
      idata_113_flg_V : in  std_logic_vector (3 downto 0);
      idata_114_flg_V : in  std_logic_vector (3 downto 0);
      idata_115_flg_V : in  std_logic_vector (3 downto 0);
      idata_116_flg_V : in  std_logic_vector (3 downto 0);
      idata_117_flg_V : in  std_logic_vector (3 downto 0);
      idata_118_flg_V : in  std_logic_vector (3 downto 0);
      idata_119_flg_V : in  std_logic_vector (3 downto 0);
      idata_120_flg_V : in  std_logic_vector (3 downto 0);
      idata_121_flg_V : in  std_logic_vector (3 downto 0);
      idata_122_flg_V : in  std_logic_vector (3 downto 0);
      idata_123_flg_V : in  std_logic_vector (3 downto 0);
      idata_124_flg_V : in  std_logic_vector (3 downto 0);
      idata_125_flg_V : in  std_logic_vector (3 downto 0);
      idata_126_flg_V : in  std_logic_vector (3 downto 0);
      idata_127_flg_V : in  std_logic_vector (3 downto 0);
      idata_128_flg_V : in  std_logic_vector (3 downto 0);
      idata_129_flg_V : in  std_logic_vector (3 downto 0);
      idata_130_flg_V : in  std_logic_vector (3 downto 0);
      idata_131_flg_V : in  std_logic_vector (3 downto 0);
      idata_132_flg_V : in  std_logic_vector (3 downto 0);
      idata_133_flg_V : in  std_logic_vector (3 downto 0);
      idata_134_flg_V : in  std_logic_vector (3 downto 0);
      idata_135_flg_V : in  std_logic_vector (3 downto 0);
      idata_136_flg_V : in  std_logic_vector (3 downto 0);
      idata_137_flg_V : in  std_logic_vector (3 downto 0);
      idata_138_flg_V : in  std_logic_vector (3 downto 0);
      idata_139_flg_V : in  std_logic_vector (3 downto 0);
      idata_140_flg_V : in  std_logic_vector (3 downto 0);
      idata_141_flg_V : in  std_logic_vector (3 downto 0);
      idata_142_flg_V : in  std_logic_vector (3 downto 0);
      idata_143_flg_V : in  std_logic_vector (3 downto 0);
      idata_144_flg_V : in  std_logic_vector (3 downto 0);
      idata_145_flg_V : in  std_logic_vector (3 downto 0);
      idata_146_flg_V : in  std_logic_vector (3 downto 0);
      idata_147_flg_V : in  std_logic_vector (3 downto 0);
      idata_148_flg_V : in  std_logic_vector (3 downto 0);
      idata_149_flg_V : in  std_logic_vector (3 downto 0);
      idata_150_flg_V : in  std_logic_vector (3 downto 0);
      idata_151_flg_V : in  std_logic_vector (3 downto 0);
      idata_152_flg_V : in  std_logic_vector (3 downto 0);
      idata_153_flg_V : in  std_logic_vector (3 downto 0);
      idata_154_flg_V : in  std_logic_vector (3 downto 0);
      idata_155_flg_V : in  std_logic_vector (3 downto 0);
      idata_156_flg_V : in  std_logic_vector (3 downto 0);
      idata_157_flg_V : in  std_logic_vector (3 downto 0);
      idata_158_flg_V : in  std_logic_vector (3 downto 0);
      idata_159_flg_V : in  std_logic_vector (3 downto 0);
      idata_160_flg_V : in  std_logic_vector (3 downto 0);
      idata_161_flg_V : in  std_logic_vector (3 downto 0);
      idata_162_flg_V : in  std_logic_vector (3 downto 0);
      idata_163_flg_V : in  std_logic_vector (3 downto 0);
      idata_164_flg_V : in  std_logic_vector (3 downto 0);
      idata_165_flg_V : in  std_logic_vector (3 downto 0);
      idata_166_flg_V : in  std_logic_vector (3 downto 0);
      idata_167_flg_V : in  std_logic_vector (3 downto 0);
      idata_168_flg_V : in  std_logic_vector (3 downto 0);
      idata_169_flg_V : in  std_logic_vector (3 downto 0);
      idata_170_flg_V : in  std_logic_vector (3 downto 0);
      idata_171_flg_V : in  std_logic_vector (3 downto 0);
      idata_172_flg_V : in  std_logic_vector (3 downto 0);
      idata_173_flg_V : in  std_logic_vector (3 downto 0);
      idata_174_flg_V : in  std_logic_vector (3 downto 0);
      idata_175_flg_V : in  std_logic_vector (3 downto 0);
      idata_176_flg_V : in  std_logic_vector (3 downto 0);
      idata_177_flg_V : in  std_logic_vector (3 downto 0);
      idata_178_flg_V : in  std_logic_vector (3 downto 0);
      idata_179_flg_V : in  std_logic_vector (3 downto 0);
      idata_180_flg_V : in  std_logic_vector (3 downto 0);
      idata_181_flg_V : in  std_logic_vector (3 downto 0);
      idata_182_flg_V : in  std_logic_vector (3 downto 0);
      idata_183_flg_V : in  std_logic_vector (3 downto 0);
      idata_184_flg_V : in  std_logic_vector (3 downto 0);
      idata_185_flg_V : in  std_logic_vector (3 downto 0);
      idata_186_flg_V : in  std_logic_vector (3 downto 0);
      idata_187_flg_V : in  std_logic_vector (3 downto 0);
      idata_188_flg_V : in  std_logic_vector (3 downto 0);
      idata_189_flg_V : in  std_logic_vector (3 downto 0);
      idata_190_flg_V : in  std_logic_vector (3 downto 0);
      idata_191_flg_V : in  std_logic_vector (3 downto 0);
      idata_192_flg_V : in  std_logic_vector (3 downto 0);
      idata_193_flg_V : in  std_logic_vector (3 downto 0);
      idata_194_flg_V : in  std_logic_vector (3 downto 0);
      idata_195_flg_V : in  std_logic_vector (3 downto 0);
      idata_196_flg_V : in  std_logic_vector (3 downto 0);
      idata_197_flg_V : in  std_logic_vector (3 downto 0);
      idata_198_flg_V : in  std_logic_vector (3 downto 0);
      idata_199_flg_V : in  std_logic_vector (3 downto 0);
      idata_200_flg_V : in  std_logic_vector (3 downto 0);
      idata_201_flg_V : in  std_logic_vector (3 downto 0);
      idata_202_flg_V : in  std_logic_vector (3 downto 0);
      idata_203_flg_V : in  std_logic_vector (3 downto 0);
      idata_204_flg_V : in  std_logic_vector (3 downto 0);
      idata_205_flg_V : in  std_logic_vector (3 downto 0);
      idata_206_flg_V : in  std_logic_vector (3 downto 0);
      idata_207_flg_V : in  std_logic_vector (3 downto 0);
      idata_208_flg_V : in  std_logic_vector (3 downto 0);
      idata_209_flg_V : in  std_logic_vector (3 downto 0);
      idata_210_flg_V : in  std_logic_vector (3 downto 0);
      idata_211_flg_V : in  std_logic_vector (3 downto 0);
      idata_212_flg_V : in  std_logic_vector (3 downto 0);
      idata_213_flg_V : in  std_logic_vector (3 downto 0);
      idata_214_flg_V : in  std_logic_vector (3 downto 0);
      idata_215_flg_V : in  std_logic_vector (3 downto 0);
      idata_216_flg_V : in  std_logic_vector (3 downto 0);
      idata_217_flg_V : in  std_logic_vector (3 downto 0);
      idata_218_flg_V : in  std_logic_vector (3 downto 0);
      idata_219_flg_V : in  std_logic_vector (3 downto 0);
      idata_220_flg_V : in  std_logic_vector (3 downto 0);
      idata_221_flg_V : in  std_logic_vector (3 downto 0);
      idata_222_flg_V : in  std_logic_vector (3 downto 0);
      idata_223_flg_V : in  std_logic_vector (3 downto 0);
      idata_224_flg_V : in  std_logic_vector (3 downto 0);
      idata_225_flg_V : in  std_logic_vector (3 downto 0);
      idata_226_flg_V : in  std_logic_vector (3 downto 0);
      idata_227_flg_V : in  std_logic_vector (3 downto 0);
      idata_228_flg_V : in  std_logic_vector (3 downto 0);
      idata_229_flg_V : in  std_logic_vector (3 downto 0);
      idata_230_flg_V : in  std_logic_vector (3 downto 0);
      idata_231_flg_V : in  std_logic_vector (3 downto 0);
      idata_232_flg_V : in  std_logic_vector (3 downto 0);
      idata_233_flg_V : in  std_logic_vector (3 downto 0);
      idata_234_flg_V : in  std_logic_vector (3 downto 0);
      idata_235_flg_V : in  std_logic_vector (3 downto 0);
      idata_236_flg_V : in  std_logic_vector (3 downto 0);
      idata_237_flg_V : in  std_logic_vector (3 downto 0);
      idata_238_flg_V : in  std_logic_vector (3 downto 0);
      idata_239_flg_V : in  std_logic_vector (3 downto 0);
      idata_240_flg_V : in  std_logic_vector (3 downto 0);
      idata_241_flg_V : in  std_logic_vector (3 downto 0);
      idata_242_flg_V : in  std_logic_vector (3 downto 0);
      idata_243_flg_V : in  std_logic_vector (3 downto 0);
      idata_244_flg_V : in  std_logic_vector (3 downto 0);
      idata_245_flg_V : in  std_logic_vector (3 downto 0);
      idata_246_flg_V : in  std_logic_vector (3 downto 0);
      idata_247_flg_V : in  std_logic_vector (3 downto 0);
      idata_248_flg_V : in  std_logic_vector (3 downto 0);
      idata_249_flg_V : in  std_logic_vector (3 downto 0);
      idata_250_flg_V : in  std_logic_vector (3 downto 0);
      idata_251_flg_V : in  std_logic_vector (3 downto 0);
      idata_252_flg_V : in  std_logic_vector (3 downto 0);
      idata_253_flg_V : in  std_logic_vector (3 downto 0);
      idata_254_flg_V : in  std_logic_vector (3 downto 0);
      idata_255_flg_V : in  std_logic_vector (3 downto 0);
      idata_256_flg_V : in  std_logic_vector (3 downto 0);
      idata_257_flg_V : in  std_logic_vector (3 downto 0);
      idata_258_flg_V : in  std_logic_vector (3 downto 0);
      idata_259_flg_V : in  std_logic_vector (3 downto 0);
      idata_260_flg_V : in  std_logic_vector (3 downto 0);
      idata_261_flg_V : in  std_logic_vector (3 downto 0);
      idata_262_flg_V : in  std_logic_vector (3 downto 0);
      idata_263_flg_V : in  std_logic_vector (3 downto 0);
      idata_264_flg_V : in  std_logic_vector (3 downto 0);
      idata_265_flg_V : in  std_logic_vector (3 downto 0);
      idata_266_flg_V : in  std_logic_vector (3 downto 0);
      idata_267_flg_V : in  std_logic_vector (3 downto 0);
      idata_268_flg_V : in  std_logic_vector (3 downto 0);
      idata_269_flg_V : in  std_logic_vector (3 downto 0);
      idata_270_flg_V : in  std_logic_vector (3 downto 0);
      idata_271_flg_V : in  std_logic_vector (3 downto 0);
      idata_272_flg_V : in  std_logic_vector (3 downto 0);
      idata_273_flg_V : in  std_logic_vector (3 downto 0);
      idata_274_flg_V : in  std_logic_vector (3 downto 0);
      idata_275_flg_V : in  std_logic_vector (3 downto 0);
      idata_276_flg_V : in  std_logic_vector (3 downto 0);
      idata_277_flg_V : in  std_logic_vector (3 downto 0);
      idata_278_flg_V : in  std_logic_vector (3 downto 0);
      idata_279_flg_V : in  std_logic_vector (3 downto 0);
      idata_280_flg_V : in  std_logic_vector (3 downto 0);
      idata_281_flg_V : in  std_logic_vector (3 downto 0);
      idata_282_flg_V : in  std_logic_vector (3 downto 0);
      idata_283_flg_V : in  std_logic_vector (3 downto 0);
      idata_284_flg_V : in  std_logic_vector (3 downto 0);
      idata_285_flg_V : in  std_logic_vector (3 downto 0);
      idata_286_flg_V : in  std_logic_vector (3 downto 0);
      idata_287_flg_V : in  std_logic_vector (3 downto 0);
      idata_288_flg_V : in  std_logic_vector (3 downto 0);
      idata_289_flg_V : in  std_logic_vector (3 downto 0);
      idata_290_flg_V : in  std_logic_vector (3 downto 0);
      idata_291_flg_V : in  std_logic_vector (3 downto 0);
      idata_292_flg_V : in  std_logic_vector (3 downto 0);
      idata_293_flg_V : in  std_logic_vector (3 downto 0);
      idata_294_flg_V : in  std_logic_vector (3 downto 0);
      idata_295_flg_V : in  std_logic_vector (3 downto 0);
      idata_296_flg_V : in  std_logic_vector (3 downto 0);
      idata_297_flg_V : in  std_logic_vector (3 downto 0);
      idata_298_flg_V : in  std_logic_vector (3 downto 0);
      idata_299_flg_V : in  std_logic_vector (3 downto 0);
      idata_300_flg_V : in  std_logic_vector (3 downto 0);
      idata_301_flg_V : in  std_logic_vector (3 downto 0);
      idata_302_flg_V : in  std_logic_vector (3 downto 0);
      idata_303_flg_V : in  std_logic_vector (3 downto 0);
      idata_304_flg_V : in  std_logic_vector (3 downto 0);
      idata_305_flg_V : in  std_logic_vector (3 downto 0);
      idata_306_flg_V : in  std_logic_vector (3 downto 0);
      idata_307_flg_V : in  std_logic_vector (3 downto 0);
      idata_308_flg_V : in  std_logic_vector (3 downto 0);
      idata_309_flg_V : in  std_logic_vector (3 downto 0);
      idata_310_flg_V : in  std_logic_vector (3 downto 0);
      idata_311_flg_V : in  std_logic_vector (3 downto 0);
      idata_312_flg_V : in  std_logic_vector (3 downto 0);
      idata_313_flg_V : in  std_logic_vector (3 downto 0);
      idata_314_flg_V : in  std_logic_vector (3 downto 0);
      idata_315_flg_V : in  std_logic_vector (3 downto 0);
      idata_316_flg_V : in  std_logic_vector (3 downto 0);
      idata_317_flg_V : in  std_logic_vector (3 downto 0);
      idata_318_flg_V : in  std_logic_vector (3 downto 0);
      idata_319_flg_V : in  std_logic_vector (3 downto 0);
      idata_320_flg_V : in  std_logic_vector (3 downto 0);
      idata_321_flg_V : in  std_logic_vector (3 downto 0);
      idata_322_flg_V : in  std_logic_vector (3 downto 0);
      idata_323_flg_V : in  std_logic_vector (3 downto 0);
      idata_324_flg_V : in  std_logic_vector (3 downto 0);
      idata_325_flg_V : in  std_logic_vector (3 downto 0);
      idata_326_flg_V : in  std_logic_vector (3 downto 0);
      idata_327_flg_V : in  std_logic_vector (3 downto 0);
      idata_328_flg_V : in  std_logic_vector (3 downto 0);
      idata_329_flg_V : in  std_logic_vector (3 downto 0);
      idata_330_flg_V : in  std_logic_vector (3 downto 0);
      idata_331_flg_V : in  std_logic_vector (3 downto 0);
      idata_332_flg_V : in  std_logic_vector (3 downto 0);
      idata_333_flg_V : in  std_logic_vector (3 downto 0);
      idata_334_flg_V : in  std_logic_vector (3 downto 0);
      idata_335_flg_V : in  std_logic_vector (3 downto 0);
      idata_336_flg_V : in  std_logic_vector (3 downto 0);
      idata_337_flg_V : in  std_logic_vector (3 downto 0);
      idata_338_flg_V : in  std_logic_vector (3 downto 0);
      idata_339_flg_V : in  std_logic_vector (3 downto 0);
      idata_340_flg_V : in  std_logic_vector (3 downto 0);
      idata_341_flg_V : in  std_logic_vector (3 downto 0);
      idata_342_flg_V : in  std_logic_vector (3 downto 0);
      idata_343_flg_V : in  std_logic_vector (3 downto 0);
      idata_344_flg_V : in  std_logic_vector (3 downto 0);
      idata_345_flg_V : in  std_logic_vector (3 downto 0);
      idata_346_flg_V : in  std_logic_vector (3 downto 0);
      idata_347_flg_V : in  std_logic_vector (3 downto 0);
      idata_348_flg_V : in  std_logic_vector (3 downto 0);
      idata_349_flg_V : in  std_logic_vector (3 downto 0);
      idata_350_flg_V : in  std_logic_vector (3 downto 0);
      idata_351_flg_V : in  std_logic_vector (3 downto 0);
      odata_0_id_V    : out std_logic_vector (8 downto 0);
      odata_1_id_V    : out std_logic_vector (8 downto 0);
      odata_2_id_V    : out std_logic_vector (8 downto 0);
      odata_3_id_V    : out std_logic_vector (8 downto 0);
      odata_4_id_V    : out std_logic_vector (8 downto 0);
      odata_5_id_V    : out std_logic_vector (8 downto 0);
      odata_6_id_V    : out std_logic_vector (8 downto 0);
      odata_7_id_V    : out std_logic_vector (8 downto 0);
      odata_8_id_V    : out std_logic_vector (8 downto 0);
      odata_9_id_V    : out std_logic_vector (8 downto 0);
      odata_10_id_V   : out std_logic_vector (8 downto 0);
      odata_11_id_V   : out std_logic_vector (8 downto 0);
      odata_12_id_V   : out std_logic_vector (8 downto 0);
      odata_13_id_V   : out std_logic_vector (8 downto 0);
      odata_14_id_V   : out std_logic_vector (8 downto 0);
      odata_15_id_V   : out std_logic_vector (8 downto 0);
      odata_0_pt_V    : out std_logic_vector (3 downto 0);
      odata_1_pt_V    : out std_logic_vector (3 downto 0);
      odata_2_pt_V    : out std_logic_vector (3 downto 0);
      odata_3_pt_V    : out std_logic_vector (3 downto 0);
      odata_4_pt_V    : out std_logic_vector (3 downto 0);
      odata_5_pt_V    : out std_logic_vector (3 downto 0);
      odata_6_pt_V    : out std_logic_vector (3 downto 0);
      odata_7_pt_V    : out std_logic_vector (3 downto 0);
      odata_8_pt_V    : out std_logic_vector (3 downto 0);
      odata_9_pt_V    : out std_logic_vector (3 downto 0);
      odata_10_pt_V   : out std_logic_vector (3 downto 0);
      odata_11_pt_V   : out std_logic_vector (3 downto 0);
      odata_12_pt_V   : out std_logic_vector (3 downto 0);
      odata_13_pt_V   : out std_logic_vector (3 downto 0);
      odata_14_pt_V   : out std_logic_vector (3 downto 0);
      odata_15_pt_V   : out std_logic_vector (3 downto 0);
      odata_0_roi_V   : out std_logic_vector (7 downto 0);
      odata_1_roi_V   : out std_logic_vector (7 downto 0);
      odata_2_roi_V   : out std_logic_vector (7 downto 0);
      odata_3_roi_V   : out std_logic_vector (7 downto 0);
      odata_4_roi_V   : out std_logic_vector (7 downto 0);
      odata_5_roi_V   : out std_logic_vector (7 downto 0);
      odata_6_roi_V   : out std_logic_vector (7 downto 0);
      odata_7_roi_V   : out std_logic_vector (7 downto 0);
      odata_8_roi_V   : out std_logic_vector (7 downto 0);
      odata_9_roi_V   : out std_logic_vector (7 downto 0);
      odata_10_roi_V  : out std_logic_vector (7 downto 0);
      odata_11_roi_V  : out std_logic_vector (7 downto 0);
      odata_12_roi_V  : out std_logic_vector (7 downto 0);
      odata_13_roi_V  : out std_logic_vector (7 downto 0);
      odata_14_roi_V  : out std_logic_vector (7 downto 0);
      odata_15_roi_V  : out std_logic_vector (7 downto 0);
      odata_0_flg_V   : out std_logic_vector (3 downto 0);
      odata_1_flg_V   : out std_logic_vector (3 downto 0);
      odata_2_flg_V   : out std_logic_vector (3 downto 0);
      odata_3_flg_V   : out std_logic_vector (3 downto 0);
      odata_4_flg_V   : out std_logic_vector (3 downto 0);
      odata_5_flg_V   : out std_logic_vector (3 downto 0);
      odata_6_flg_V   : out std_logic_vector (3 downto 0);
      odata_7_flg_V   : out std_logic_vector (3 downto 0);
      odata_8_flg_V   : out std_logic_vector (3 downto 0);
      odata_9_flg_V   : out std_logic_vector (3 downto 0);
      odata_10_flg_V  : out std_logic_vector (3 downto 0);
      odata_11_flg_V  : out std_logic_vector (3 downto 0);
      odata_12_flg_V  : out std_logic_vector (3 downto 0);
      odata_13_flg_V  : out std_logic_vector (3 downto 0);
      odata_14_flg_V  : out std_logic_vector (3 downto 0);
      odata_15_flg_V  : out std_logic_vector (3 downto 0));
  end component compare_main;

  -- registered signals


  signal ap_start_reg : std_logic;

  signal idata_0_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_1_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_2_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_3_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_4_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_5_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_6_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_7_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_8_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_9_pt_V_reg    : std_logic_vector (3 downto 0);
  signal idata_10_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_11_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_12_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_13_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_14_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_15_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_16_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_17_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_18_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_19_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_20_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_21_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_22_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_23_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_24_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_25_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_26_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_27_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_28_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_29_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_30_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_31_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_32_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_33_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_34_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_35_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_36_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_37_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_38_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_39_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_40_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_41_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_42_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_43_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_44_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_45_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_46_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_47_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_48_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_49_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_50_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_51_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_52_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_53_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_54_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_55_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_56_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_57_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_58_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_59_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_60_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_61_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_62_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_63_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_64_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_65_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_66_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_67_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_68_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_69_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_70_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_71_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_72_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_73_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_74_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_75_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_76_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_77_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_78_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_79_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_80_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_81_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_82_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_83_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_84_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_85_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_86_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_87_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_88_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_89_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_90_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_91_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_92_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_93_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_94_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_95_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_96_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_97_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_98_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_99_pt_V_reg   : std_logic_vector (3 downto 0);
  signal idata_100_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_101_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_102_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_103_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_104_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_105_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_106_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_107_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_108_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_109_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_110_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_111_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_112_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_113_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_114_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_115_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_116_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_117_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_118_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_119_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_120_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_121_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_122_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_123_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_124_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_125_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_126_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_127_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_128_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_129_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_130_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_131_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_132_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_133_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_134_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_135_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_136_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_137_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_138_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_139_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_140_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_141_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_142_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_143_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_144_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_145_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_146_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_147_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_148_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_149_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_150_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_151_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_152_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_153_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_154_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_155_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_156_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_157_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_158_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_159_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_160_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_161_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_162_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_163_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_164_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_165_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_166_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_167_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_168_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_169_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_170_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_171_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_172_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_173_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_174_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_175_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_176_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_177_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_178_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_179_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_180_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_181_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_182_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_183_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_184_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_185_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_186_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_187_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_188_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_189_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_190_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_191_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_192_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_193_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_194_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_195_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_196_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_197_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_198_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_199_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_200_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_201_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_202_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_203_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_204_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_205_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_206_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_207_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_208_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_209_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_210_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_211_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_212_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_213_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_214_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_215_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_216_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_217_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_218_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_219_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_220_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_221_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_222_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_223_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_224_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_225_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_226_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_227_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_228_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_229_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_230_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_231_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_232_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_233_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_234_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_235_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_236_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_237_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_238_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_239_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_240_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_241_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_242_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_243_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_244_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_245_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_246_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_247_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_248_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_249_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_250_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_251_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_252_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_253_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_254_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_255_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_256_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_257_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_258_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_259_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_260_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_261_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_262_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_263_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_264_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_265_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_266_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_267_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_268_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_269_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_270_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_271_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_272_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_273_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_274_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_275_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_276_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_277_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_278_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_279_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_280_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_281_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_282_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_283_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_284_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_285_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_286_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_287_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_288_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_289_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_290_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_291_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_292_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_293_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_294_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_295_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_296_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_297_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_298_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_299_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_300_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_301_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_302_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_303_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_304_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_305_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_306_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_307_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_308_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_309_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_310_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_311_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_312_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_313_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_314_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_315_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_316_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_317_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_318_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_319_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_320_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_321_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_322_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_323_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_324_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_325_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_326_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_327_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_328_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_329_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_330_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_331_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_332_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_333_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_334_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_335_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_336_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_337_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_338_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_339_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_340_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_341_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_342_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_343_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_344_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_345_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_346_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_347_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_348_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_349_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_350_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_351_pt_V_reg  : std_logic_vector (3 downto 0);
  signal idata_0_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_1_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_2_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_3_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_4_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_5_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_6_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_7_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_8_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_9_roi_V_reg   : std_logic_vector (7 downto 0);
  signal idata_10_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_11_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_12_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_13_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_14_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_15_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_16_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_17_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_18_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_19_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_20_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_21_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_22_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_23_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_24_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_25_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_26_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_27_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_28_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_29_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_30_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_31_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_32_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_33_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_34_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_35_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_36_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_37_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_38_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_39_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_40_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_41_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_42_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_43_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_44_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_45_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_46_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_47_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_48_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_49_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_50_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_51_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_52_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_53_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_54_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_55_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_56_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_57_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_58_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_59_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_60_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_61_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_62_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_63_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_64_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_65_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_66_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_67_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_68_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_69_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_70_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_71_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_72_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_73_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_74_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_75_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_76_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_77_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_78_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_79_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_80_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_81_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_82_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_83_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_84_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_85_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_86_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_87_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_88_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_89_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_90_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_91_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_92_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_93_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_94_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_95_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_96_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_97_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_98_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_99_roi_V_reg  : std_logic_vector (7 downto 0);
  signal idata_100_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_101_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_102_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_103_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_104_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_105_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_106_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_107_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_108_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_109_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_110_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_111_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_112_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_113_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_114_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_115_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_116_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_117_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_118_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_119_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_120_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_121_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_122_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_123_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_124_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_125_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_126_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_127_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_128_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_129_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_130_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_131_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_132_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_133_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_134_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_135_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_136_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_137_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_138_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_139_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_140_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_141_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_142_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_143_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_144_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_145_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_146_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_147_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_148_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_149_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_150_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_151_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_152_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_153_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_154_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_155_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_156_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_157_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_158_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_159_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_160_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_161_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_162_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_163_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_164_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_165_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_166_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_167_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_168_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_169_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_170_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_171_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_172_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_173_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_174_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_175_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_176_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_177_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_178_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_179_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_180_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_181_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_182_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_183_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_184_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_185_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_186_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_187_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_188_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_189_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_190_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_191_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_192_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_193_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_194_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_195_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_196_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_197_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_198_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_199_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_200_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_201_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_202_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_203_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_204_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_205_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_206_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_207_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_208_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_209_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_210_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_211_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_212_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_213_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_214_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_215_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_216_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_217_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_218_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_219_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_220_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_221_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_222_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_223_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_224_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_225_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_226_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_227_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_228_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_229_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_230_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_231_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_232_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_233_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_234_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_235_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_236_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_237_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_238_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_239_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_240_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_241_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_242_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_243_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_244_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_245_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_246_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_247_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_248_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_249_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_250_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_251_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_252_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_253_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_254_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_255_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_256_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_257_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_258_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_259_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_260_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_261_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_262_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_263_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_264_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_265_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_266_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_267_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_268_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_269_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_270_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_271_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_272_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_273_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_274_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_275_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_276_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_277_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_278_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_279_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_280_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_281_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_282_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_283_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_284_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_285_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_286_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_287_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_288_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_289_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_290_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_291_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_292_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_293_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_294_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_295_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_296_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_297_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_298_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_299_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_300_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_301_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_302_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_303_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_304_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_305_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_306_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_307_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_308_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_309_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_310_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_311_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_312_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_313_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_314_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_315_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_316_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_317_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_318_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_319_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_320_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_321_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_322_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_323_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_324_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_325_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_326_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_327_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_328_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_329_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_330_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_331_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_332_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_333_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_334_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_335_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_336_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_337_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_338_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_339_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_340_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_341_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_342_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_343_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_344_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_345_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_346_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_347_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_348_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_349_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_350_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_351_roi_V_reg : std_logic_vector (7 downto 0);
  signal idata_0_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_1_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_2_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_3_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_4_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_5_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_6_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_7_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_8_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_9_flg_V_reg   : std_logic_vector (3 downto 0);
  signal idata_10_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_11_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_12_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_13_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_14_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_15_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_16_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_17_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_18_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_19_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_20_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_21_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_22_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_23_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_24_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_25_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_26_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_27_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_28_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_29_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_30_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_31_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_32_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_33_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_34_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_35_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_36_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_37_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_38_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_39_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_40_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_41_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_42_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_43_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_44_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_45_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_46_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_47_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_48_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_49_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_50_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_51_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_52_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_53_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_54_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_55_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_56_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_57_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_58_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_59_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_60_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_61_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_62_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_63_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_64_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_65_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_66_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_67_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_68_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_69_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_70_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_71_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_72_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_73_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_74_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_75_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_76_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_77_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_78_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_79_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_80_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_81_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_82_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_83_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_84_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_85_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_86_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_87_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_88_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_89_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_90_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_91_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_92_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_93_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_94_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_95_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_96_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_97_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_98_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_99_flg_V_reg  : std_logic_vector (3 downto 0);
  signal idata_100_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_101_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_102_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_103_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_104_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_105_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_106_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_107_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_108_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_109_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_110_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_111_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_112_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_113_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_114_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_115_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_116_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_117_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_118_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_119_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_120_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_121_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_122_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_123_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_124_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_125_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_126_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_127_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_128_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_129_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_130_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_131_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_132_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_133_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_134_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_135_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_136_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_137_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_138_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_139_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_140_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_141_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_142_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_143_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_144_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_145_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_146_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_147_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_148_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_149_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_150_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_151_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_152_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_153_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_154_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_155_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_156_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_157_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_158_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_159_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_160_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_161_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_162_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_163_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_164_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_165_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_166_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_167_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_168_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_169_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_170_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_171_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_172_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_173_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_174_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_175_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_176_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_177_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_178_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_179_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_180_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_181_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_182_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_183_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_184_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_185_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_186_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_187_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_188_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_189_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_190_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_191_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_192_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_193_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_194_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_195_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_196_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_197_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_198_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_199_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_200_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_201_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_202_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_203_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_204_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_205_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_206_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_207_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_208_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_209_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_210_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_211_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_212_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_213_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_214_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_215_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_216_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_217_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_218_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_219_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_220_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_221_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_222_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_223_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_224_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_225_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_226_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_227_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_228_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_229_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_230_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_231_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_232_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_233_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_234_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_235_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_236_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_237_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_238_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_239_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_240_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_241_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_242_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_243_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_244_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_245_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_246_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_247_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_248_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_249_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_250_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_251_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_252_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_253_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_254_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_255_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_256_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_257_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_258_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_259_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_260_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_261_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_262_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_263_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_264_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_265_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_266_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_267_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_268_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_269_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_270_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_271_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_272_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_273_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_274_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_275_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_276_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_277_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_278_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_279_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_280_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_281_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_282_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_283_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_284_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_285_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_286_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_287_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_288_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_289_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_290_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_291_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_292_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_293_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_294_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_295_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_296_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_297_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_298_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_299_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_300_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_301_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_302_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_303_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_304_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_305_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_306_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_307_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_308_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_309_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_310_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_311_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_312_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_313_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_314_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_315_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_316_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_317_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_318_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_319_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_320_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_321_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_322_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_323_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_324_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_325_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_326_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_327_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_328_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_329_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_330_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_331_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_332_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_333_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_334_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_335_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_336_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_337_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_338_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_339_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_340_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_341_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_342_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_343_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_344_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_345_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_346_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_347_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_348_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_349_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_350_flg_V_reg : std_logic_vector (3 downto 0);
  signal idata_351_flg_V_reg : std_logic_vector (3 downto 0);


begin  -- architecture rtl

  --in reg
  reg_p : process (ap_clk) is
  begin
    if rising_edge(ap_clk) then

      ap_start_reg        <= ap_start;
      idata_0_pt_V_reg    <= idata_0_pt_V;
      idata_1_pt_V_reg    <= idata_1_pt_V;
      idata_2_pt_V_reg    <= idata_2_pt_V;
      idata_3_pt_V_reg    <= idata_3_pt_V;
      idata_4_pt_V_reg    <= idata_4_pt_V;
      idata_5_pt_V_reg    <= idata_5_pt_V;
      idata_6_pt_V_reg    <= idata_6_pt_V;
      idata_7_pt_V_reg    <= idata_7_pt_V;
      idata_8_pt_V_reg    <= idata_8_pt_V;
      idata_9_pt_V_reg    <= idata_9_pt_V;
      idata_10_pt_V_reg   <= idata_10_pt_V;
      idata_11_pt_V_reg   <= idata_11_pt_V;
      idata_12_pt_V_reg   <= idata_12_pt_V;
      idata_13_pt_V_reg   <= idata_13_pt_V;
      idata_14_pt_V_reg   <= idata_14_pt_V;
      idata_15_pt_V_reg   <= idata_15_pt_V;
      idata_16_pt_V_reg   <= idata_16_pt_V;
      idata_17_pt_V_reg   <= idata_17_pt_V;
      idata_18_pt_V_reg   <= idata_18_pt_V;
      idata_19_pt_V_reg   <= idata_19_pt_V;
      idata_20_pt_V_reg   <= idata_20_pt_V;
      idata_21_pt_V_reg   <= idata_21_pt_V;
      idata_22_pt_V_reg   <= idata_22_pt_V;
      idata_23_pt_V_reg   <= idata_23_pt_V;
      idata_24_pt_V_reg   <= idata_24_pt_V;
      idata_25_pt_V_reg   <= idata_25_pt_V;
      idata_26_pt_V_reg   <= idata_26_pt_V;
      idata_27_pt_V_reg   <= idata_27_pt_V;
      idata_28_pt_V_reg   <= idata_28_pt_V;
      idata_29_pt_V_reg   <= idata_29_pt_V;
      idata_30_pt_V_reg   <= idata_30_pt_V;
      idata_31_pt_V_reg   <= idata_31_pt_V;
      idata_32_pt_V_reg   <= idata_32_pt_V;
      idata_33_pt_V_reg   <= idata_33_pt_V;
      idata_34_pt_V_reg   <= idata_34_pt_V;
      idata_35_pt_V_reg   <= idata_35_pt_V;
      idata_36_pt_V_reg   <= idata_36_pt_V;
      idata_37_pt_V_reg   <= idata_37_pt_V;
      idata_38_pt_V_reg   <= idata_38_pt_V;
      idata_39_pt_V_reg   <= idata_39_pt_V;
      idata_40_pt_V_reg   <= idata_40_pt_V;
      idata_41_pt_V_reg   <= idata_41_pt_V;
      idata_42_pt_V_reg   <= idata_42_pt_V;
      idata_43_pt_V_reg   <= idata_43_pt_V;
      idata_44_pt_V_reg   <= idata_44_pt_V;
      idata_45_pt_V_reg   <= idata_45_pt_V;
      idata_46_pt_V_reg   <= idata_46_pt_V;
      idata_47_pt_V_reg   <= idata_47_pt_V;
      idata_48_pt_V_reg   <= idata_48_pt_V;
      idata_49_pt_V_reg   <= idata_49_pt_V;
      idata_50_pt_V_reg   <= idata_50_pt_V;
      idata_51_pt_V_reg   <= idata_51_pt_V;
      idata_52_pt_V_reg   <= idata_52_pt_V;
      idata_53_pt_V_reg   <= idata_53_pt_V;
      idata_54_pt_V_reg   <= idata_54_pt_V;
      idata_55_pt_V_reg   <= idata_55_pt_V;
      idata_56_pt_V_reg   <= idata_56_pt_V;
      idata_57_pt_V_reg   <= idata_57_pt_V;
      idata_58_pt_V_reg   <= idata_58_pt_V;
      idata_59_pt_V_reg   <= idata_59_pt_V;
      idata_60_pt_V_reg   <= idata_60_pt_V;
      idata_61_pt_V_reg   <= idata_61_pt_V;
      idata_62_pt_V_reg   <= idata_62_pt_V;
      idata_63_pt_V_reg   <= idata_63_pt_V;
      idata_64_pt_V_reg   <= idata_64_pt_V;
      idata_65_pt_V_reg   <= idata_65_pt_V;
      idata_66_pt_V_reg   <= idata_66_pt_V;
      idata_67_pt_V_reg   <= idata_67_pt_V;
      idata_68_pt_V_reg   <= idata_68_pt_V;
      idata_69_pt_V_reg   <= idata_69_pt_V;
      idata_70_pt_V_reg   <= idata_70_pt_V;
      idata_71_pt_V_reg   <= idata_71_pt_V;
      idata_72_pt_V_reg   <= idata_72_pt_V;
      idata_73_pt_V_reg   <= idata_73_pt_V;
      idata_74_pt_V_reg   <= idata_74_pt_V;
      idata_75_pt_V_reg   <= idata_75_pt_V;
      idata_76_pt_V_reg   <= idata_76_pt_V;
      idata_77_pt_V_reg   <= idata_77_pt_V;
      idata_78_pt_V_reg   <= idata_78_pt_V;
      idata_79_pt_V_reg   <= idata_79_pt_V;
      idata_80_pt_V_reg   <= idata_80_pt_V;
      idata_81_pt_V_reg   <= idata_81_pt_V;
      idata_82_pt_V_reg   <= idata_82_pt_V;
      idata_83_pt_V_reg   <= idata_83_pt_V;
      idata_84_pt_V_reg   <= idata_84_pt_V;
      idata_85_pt_V_reg   <= idata_85_pt_V;
      idata_86_pt_V_reg   <= idata_86_pt_V;
      idata_87_pt_V_reg   <= idata_87_pt_V;
      idata_88_pt_V_reg   <= idata_88_pt_V;
      idata_89_pt_V_reg   <= idata_89_pt_V;
      idata_90_pt_V_reg   <= idata_90_pt_V;
      idata_91_pt_V_reg   <= idata_91_pt_V;
      idata_92_pt_V_reg   <= idata_92_pt_V;
      idata_93_pt_V_reg   <= idata_93_pt_V;
      idata_94_pt_V_reg   <= idata_94_pt_V;
      idata_95_pt_V_reg   <= idata_95_pt_V;
      idata_96_pt_V_reg   <= idata_96_pt_V;
      idata_97_pt_V_reg   <= idata_97_pt_V;
      idata_98_pt_V_reg   <= idata_98_pt_V;
      idata_99_pt_V_reg   <= idata_99_pt_V;
      idata_100_pt_V_reg  <= idata_100_pt_V;
      idata_101_pt_V_reg  <= idata_101_pt_V;
      idata_102_pt_V_reg  <= idata_102_pt_V;
      idata_103_pt_V_reg  <= idata_103_pt_V;
      idata_104_pt_V_reg  <= idata_104_pt_V;
      idata_105_pt_V_reg  <= idata_105_pt_V;
      idata_106_pt_V_reg  <= idata_106_pt_V;
      idata_107_pt_V_reg  <= idata_107_pt_V;
      idata_108_pt_V_reg  <= idata_108_pt_V;
      idata_109_pt_V_reg  <= idata_109_pt_V;
      idata_110_pt_V_reg  <= idata_110_pt_V;
      idata_111_pt_V_reg  <= idata_111_pt_V;
      idata_112_pt_V_reg  <= idata_112_pt_V;
      idata_113_pt_V_reg  <= idata_113_pt_V;
      idata_114_pt_V_reg  <= idata_114_pt_V;
      idata_115_pt_V_reg  <= idata_115_pt_V;
      idata_116_pt_V_reg  <= idata_116_pt_V;
      idata_117_pt_V_reg  <= idata_117_pt_V;
      idata_118_pt_V_reg  <= idata_118_pt_V;
      idata_119_pt_V_reg  <= idata_119_pt_V;
      idata_120_pt_V_reg  <= idata_120_pt_V;
      idata_121_pt_V_reg  <= idata_121_pt_V;
      idata_122_pt_V_reg  <= idata_122_pt_V;
      idata_123_pt_V_reg  <= idata_123_pt_V;
      idata_124_pt_V_reg  <= idata_124_pt_V;
      idata_125_pt_V_reg  <= idata_125_pt_V;
      idata_126_pt_V_reg  <= idata_126_pt_V;
      idata_127_pt_V_reg  <= idata_127_pt_V;
      idata_128_pt_V_reg  <= idata_128_pt_V;
      idata_129_pt_V_reg  <= idata_129_pt_V;
      idata_130_pt_V_reg  <= idata_130_pt_V;
      idata_131_pt_V_reg  <= idata_131_pt_V;
      idata_132_pt_V_reg  <= idata_132_pt_V;
      idata_133_pt_V_reg  <= idata_133_pt_V;
      idata_134_pt_V_reg  <= idata_134_pt_V;
      idata_135_pt_V_reg  <= idata_135_pt_V;
      idata_136_pt_V_reg  <= idata_136_pt_V;
      idata_137_pt_V_reg  <= idata_137_pt_V;
      idata_138_pt_V_reg  <= idata_138_pt_V;
      idata_139_pt_V_reg  <= idata_139_pt_V;
      idata_140_pt_V_reg  <= idata_140_pt_V;
      idata_141_pt_V_reg  <= idata_141_pt_V;
      idata_142_pt_V_reg  <= idata_142_pt_V;
      idata_143_pt_V_reg  <= idata_143_pt_V;
      idata_144_pt_V_reg  <= idata_144_pt_V;
      idata_145_pt_V_reg  <= idata_145_pt_V;
      idata_146_pt_V_reg  <= idata_146_pt_V;
      idata_147_pt_V_reg  <= idata_147_pt_V;
      idata_148_pt_V_reg  <= idata_148_pt_V;
      idata_149_pt_V_reg  <= idata_149_pt_V;
      idata_150_pt_V_reg  <= idata_150_pt_V;
      idata_151_pt_V_reg  <= idata_151_pt_V;
      idata_152_pt_V_reg  <= idata_152_pt_V;
      idata_153_pt_V_reg  <= idata_153_pt_V;
      idata_154_pt_V_reg  <= idata_154_pt_V;
      idata_155_pt_V_reg  <= idata_155_pt_V;
      idata_156_pt_V_reg  <= idata_156_pt_V;
      idata_157_pt_V_reg  <= idata_157_pt_V;
      idata_158_pt_V_reg  <= idata_158_pt_V;
      idata_159_pt_V_reg  <= idata_159_pt_V;
      idata_160_pt_V_reg  <= idata_160_pt_V;
      idata_161_pt_V_reg  <= idata_161_pt_V;
      idata_162_pt_V_reg  <= idata_162_pt_V;
      idata_163_pt_V_reg  <= idata_163_pt_V;
      idata_164_pt_V_reg  <= idata_164_pt_V;
      idata_165_pt_V_reg  <= idata_165_pt_V;
      idata_166_pt_V_reg  <= idata_166_pt_V;
      idata_167_pt_V_reg  <= idata_167_pt_V;
      idata_168_pt_V_reg  <= idata_168_pt_V;
      idata_169_pt_V_reg  <= idata_169_pt_V;
      idata_170_pt_V_reg  <= idata_170_pt_V;
      idata_171_pt_V_reg  <= idata_171_pt_V;
      idata_172_pt_V_reg  <= idata_172_pt_V;
      idata_173_pt_V_reg  <= idata_173_pt_V;
      idata_174_pt_V_reg  <= idata_174_pt_V;
      idata_175_pt_V_reg  <= idata_175_pt_V;
      idata_176_pt_V_reg  <= idata_176_pt_V;
      idata_177_pt_V_reg  <= idata_177_pt_V;
      idata_178_pt_V_reg  <= idata_178_pt_V;
      idata_179_pt_V_reg  <= idata_179_pt_V;
      idata_180_pt_V_reg  <= idata_180_pt_V;
      idata_181_pt_V_reg  <= idata_181_pt_V;
      idata_182_pt_V_reg  <= idata_182_pt_V;
      idata_183_pt_V_reg  <= idata_183_pt_V;
      idata_184_pt_V_reg  <= idata_184_pt_V;
      idata_185_pt_V_reg  <= idata_185_pt_V;
      idata_186_pt_V_reg  <= idata_186_pt_V;
      idata_187_pt_V_reg  <= idata_187_pt_V;
      idata_188_pt_V_reg  <= idata_188_pt_V;
      idata_189_pt_V_reg  <= idata_189_pt_V;
      idata_190_pt_V_reg  <= idata_190_pt_V;
      idata_191_pt_V_reg  <= idata_191_pt_V;
      idata_192_pt_V_reg  <= idata_192_pt_V;
      idata_193_pt_V_reg  <= idata_193_pt_V;
      idata_194_pt_V_reg  <= idata_194_pt_V;
      idata_195_pt_V_reg  <= idata_195_pt_V;
      idata_196_pt_V_reg  <= idata_196_pt_V;
      idata_197_pt_V_reg  <= idata_197_pt_V;
      idata_198_pt_V_reg  <= idata_198_pt_V;
      idata_199_pt_V_reg  <= idata_199_pt_V;
      idata_200_pt_V_reg  <= idata_200_pt_V;
      idata_201_pt_V_reg  <= idata_201_pt_V;
      idata_202_pt_V_reg  <= idata_202_pt_V;
      idata_203_pt_V_reg  <= idata_203_pt_V;
      idata_204_pt_V_reg  <= idata_204_pt_V;
      idata_205_pt_V_reg  <= idata_205_pt_V;
      idata_206_pt_V_reg  <= idata_206_pt_V;
      idata_207_pt_V_reg  <= idata_207_pt_V;
      idata_208_pt_V_reg  <= idata_208_pt_V;
      idata_209_pt_V_reg  <= idata_209_pt_V;
      idata_210_pt_V_reg  <= idata_210_pt_V;
      idata_211_pt_V_reg  <= idata_211_pt_V;
      idata_212_pt_V_reg  <= idata_212_pt_V;
      idata_213_pt_V_reg  <= idata_213_pt_V;
      idata_214_pt_V_reg  <= idata_214_pt_V;
      idata_215_pt_V_reg  <= idata_215_pt_V;
      idata_216_pt_V_reg  <= idata_216_pt_V;
      idata_217_pt_V_reg  <= idata_217_pt_V;
      idata_218_pt_V_reg  <= idata_218_pt_V;
      idata_219_pt_V_reg  <= idata_219_pt_V;
      idata_220_pt_V_reg  <= idata_220_pt_V;
      idata_221_pt_V_reg  <= idata_221_pt_V;
      idata_222_pt_V_reg  <= idata_222_pt_V;
      idata_223_pt_V_reg  <= idata_223_pt_V;
      idata_224_pt_V_reg  <= idata_224_pt_V;
      idata_225_pt_V_reg  <= idata_225_pt_V;
      idata_226_pt_V_reg  <= idata_226_pt_V;
      idata_227_pt_V_reg  <= idata_227_pt_V;
      idata_228_pt_V_reg  <= idata_228_pt_V;
      idata_229_pt_V_reg  <= idata_229_pt_V;
      idata_230_pt_V_reg  <= idata_230_pt_V;
      idata_231_pt_V_reg  <= idata_231_pt_V;
      idata_232_pt_V_reg  <= idata_232_pt_V;
      idata_233_pt_V_reg  <= idata_233_pt_V;
      idata_234_pt_V_reg  <= idata_234_pt_V;
      idata_235_pt_V_reg  <= idata_235_pt_V;
      idata_236_pt_V_reg  <= idata_236_pt_V;
      idata_237_pt_V_reg  <= idata_237_pt_V;
      idata_238_pt_V_reg  <= idata_238_pt_V;
      idata_239_pt_V_reg  <= idata_239_pt_V;
      idata_240_pt_V_reg  <= idata_240_pt_V;
      idata_241_pt_V_reg  <= idata_241_pt_V;
      idata_242_pt_V_reg  <= idata_242_pt_V;
      idata_243_pt_V_reg  <= idata_243_pt_V;
      idata_244_pt_V_reg  <= idata_244_pt_V;
      idata_245_pt_V_reg  <= idata_245_pt_V;
      idata_246_pt_V_reg  <= idata_246_pt_V;
      idata_247_pt_V_reg  <= idata_247_pt_V;
      idata_248_pt_V_reg  <= idata_248_pt_V;
      idata_249_pt_V_reg  <= idata_249_pt_V;
      idata_250_pt_V_reg  <= idata_250_pt_V;
      idata_251_pt_V_reg  <= idata_251_pt_V;
      idata_252_pt_V_reg  <= idata_252_pt_V;
      idata_253_pt_V_reg  <= idata_253_pt_V;
      idata_254_pt_V_reg  <= idata_254_pt_V;
      idata_255_pt_V_reg  <= idata_255_pt_V;
      idata_256_pt_V_reg  <= idata_256_pt_V;
      idata_257_pt_V_reg  <= idata_257_pt_V;
      idata_258_pt_V_reg  <= idata_258_pt_V;
      idata_259_pt_V_reg  <= idata_259_pt_V;
      idata_260_pt_V_reg  <= idata_260_pt_V;
      idata_261_pt_V_reg  <= idata_261_pt_V;
      idata_262_pt_V_reg  <= idata_262_pt_V;
      idata_263_pt_V_reg  <= idata_263_pt_V;
      idata_264_pt_V_reg  <= idata_264_pt_V;
      idata_265_pt_V_reg  <= idata_265_pt_V;
      idata_266_pt_V_reg  <= idata_266_pt_V;
      idata_267_pt_V_reg  <= idata_267_pt_V;
      idata_268_pt_V_reg  <= idata_268_pt_V;
      idata_269_pt_V_reg  <= idata_269_pt_V;
      idata_270_pt_V_reg  <= idata_270_pt_V;
      idata_271_pt_V_reg  <= idata_271_pt_V;
      idata_272_pt_V_reg  <= idata_272_pt_V;
      idata_273_pt_V_reg  <= idata_273_pt_V;
      idata_274_pt_V_reg  <= idata_274_pt_V;
      idata_275_pt_V_reg  <= idata_275_pt_V;
      idata_276_pt_V_reg  <= idata_276_pt_V;
      idata_277_pt_V_reg  <= idata_277_pt_V;
      idata_278_pt_V_reg  <= idata_278_pt_V;
      idata_279_pt_V_reg  <= idata_279_pt_V;
      idata_280_pt_V_reg  <= idata_280_pt_V;
      idata_281_pt_V_reg  <= idata_281_pt_V;
      idata_282_pt_V_reg  <= idata_282_pt_V;
      idata_283_pt_V_reg  <= idata_283_pt_V;
      idata_284_pt_V_reg  <= idata_284_pt_V;
      idata_285_pt_V_reg  <= idata_285_pt_V;
      idata_286_pt_V_reg  <= idata_286_pt_V;
      idata_287_pt_V_reg  <= idata_287_pt_V;
      idata_288_pt_V_reg  <= idata_288_pt_V;
      idata_289_pt_V_reg  <= idata_289_pt_V;
      idata_290_pt_V_reg  <= idata_290_pt_V;
      idata_291_pt_V_reg  <= idata_291_pt_V;
      idata_292_pt_V_reg  <= idata_292_pt_V;
      idata_293_pt_V_reg  <= idata_293_pt_V;
      idata_294_pt_V_reg  <= idata_294_pt_V;
      idata_295_pt_V_reg  <= idata_295_pt_V;
      idata_296_pt_V_reg  <= idata_296_pt_V;
      idata_297_pt_V_reg  <= idata_297_pt_V;
      idata_298_pt_V_reg  <= idata_298_pt_V;
      idata_299_pt_V_reg  <= idata_299_pt_V;
      idata_300_pt_V_reg  <= idata_300_pt_V;
      idata_301_pt_V_reg  <= idata_301_pt_V;
      idata_302_pt_V_reg  <= idata_302_pt_V;
      idata_303_pt_V_reg  <= idata_303_pt_V;
      idata_304_pt_V_reg  <= idata_304_pt_V;
      idata_305_pt_V_reg  <= idata_305_pt_V;
      idata_306_pt_V_reg  <= idata_306_pt_V;
      idata_307_pt_V_reg  <= idata_307_pt_V;
      idata_308_pt_V_reg  <= idata_308_pt_V;
      idata_309_pt_V_reg  <= idata_309_pt_V;
      idata_310_pt_V_reg  <= idata_310_pt_V;
      idata_311_pt_V_reg  <= idata_311_pt_V;
      idata_312_pt_V_reg  <= idata_312_pt_V;
      idata_313_pt_V_reg  <= idata_313_pt_V;
      idata_314_pt_V_reg  <= idata_314_pt_V;
      idata_315_pt_V_reg  <= idata_315_pt_V;
      idata_316_pt_V_reg  <= idata_316_pt_V;
      idata_317_pt_V_reg  <= idata_317_pt_V;
      idata_318_pt_V_reg  <= idata_318_pt_V;
      idata_319_pt_V_reg  <= idata_319_pt_V;
      idata_320_pt_V_reg  <= idata_320_pt_V;
      idata_321_pt_V_reg  <= idata_321_pt_V;
      idata_322_pt_V_reg  <= idata_322_pt_V;
      idata_323_pt_V_reg  <= idata_323_pt_V;
      idata_324_pt_V_reg  <= idata_324_pt_V;
      idata_325_pt_V_reg  <= idata_325_pt_V;
      idata_326_pt_V_reg  <= idata_326_pt_V;
      idata_327_pt_V_reg  <= idata_327_pt_V;
      idata_328_pt_V_reg  <= idata_328_pt_V;
      idata_329_pt_V_reg  <= idata_329_pt_V;
      idata_330_pt_V_reg  <= idata_330_pt_V;
      idata_331_pt_V_reg  <= idata_331_pt_V;
      idata_332_pt_V_reg  <= idata_332_pt_V;
      idata_333_pt_V_reg  <= idata_333_pt_V;
      idata_334_pt_V_reg  <= idata_334_pt_V;
      idata_335_pt_V_reg  <= idata_335_pt_V;
      idata_336_pt_V_reg  <= idata_336_pt_V;
      idata_337_pt_V_reg  <= idata_337_pt_V;
      idata_338_pt_V_reg  <= idata_338_pt_V;
      idata_339_pt_V_reg  <= idata_339_pt_V;
      idata_340_pt_V_reg  <= idata_340_pt_V;
      idata_341_pt_V_reg  <= idata_341_pt_V;
      idata_342_pt_V_reg  <= idata_342_pt_V;
      idata_343_pt_V_reg  <= idata_343_pt_V;
      idata_344_pt_V_reg  <= idata_344_pt_V;
      idata_345_pt_V_reg  <= idata_345_pt_V;
      idata_346_pt_V_reg  <= idata_346_pt_V;
      idata_347_pt_V_reg  <= idata_347_pt_V;
      idata_348_pt_V_reg  <= idata_348_pt_V;
      idata_349_pt_V_reg  <= idata_349_pt_V;
      idata_350_pt_V_reg  <= idata_350_pt_V;
      idata_351_pt_V_reg  <= idata_351_pt_V;
      idata_0_roi_V_reg   <= idata_0_roi_V;
      idata_1_roi_V_reg   <= idata_1_roi_V;
      idata_2_roi_V_reg   <= idata_2_roi_V;
      idata_3_roi_V_reg   <= idata_3_roi_V;
      idata_4_roi_V_reg   <= idata_4_roi_V;
      idata_5_roi_V_reg   <= idata_5_roi_V;
      idata_6_roi_V_reg   <= idata_6_roi_V;
      idata_7_roi_V_reg   <= idata_7_roi_V;
      idata_8_roi_V_reg   <= idata_8_roi_V;
      idata_9_roi_V_reg   <= idata_9_roi_V;
      idata_10_roi_V_reg  <= idata_10_roi_V;
      idata_11_roi_V_reg  <= idata_11_roi_V;
      idata_12_roi_V_reg  <= idata_12_roi_V;
      idata_13_roi_V_reg  <= idata_13_roi_V;
      idata_14_roi_V_reg  <= idata_14_roi_V;
      idata_15_roi_V_reg  <= idata_15_roi_V;
      idata_16_roi_V_reg  <= idata_16_roi_V;
      idata_17_roi_V_reg  <= idata_17_roi_V;
      idata_18_roi_V_reg  <= idata_18_roi_V;
      idata_19_roi_V_reg  <= idata_19_roi_V;
      idata_20_roi_V_reg  <= idata_20_roi_V;
      idata_21_roi_V_reg  <= idata_21_roi_V;
      idata_22_roi_V_reg  <= idata_22_roi_V;
      idata_23_roi_V_reg  <= idata_23_roi_V;
      idata_24_roi_V_reg  <= idata_24_roi_V;
      idata_25_roi_V_reg  <= idata_25_roi_V;
      idata_26_roi_V_reg  <= idata_26_roi_V;
      idata_27_roi_V_reg  <= idata_27_roi_V;
      idata_28_roi_V_reg  <= idata_28_roi_V;
      idata_29_roi_V_reg  <= idata_29_roi_V;
      idata_30_roi_V_reg  <= idata_30_roi_V;
      idata_31_roi_V_reg  <= idata_31_roi_V;
      idata_32_roi_V_reg  <= idata_32_roi_V;
      idata_33_roi_V_reg  <= idata_33_roi_V;
      idata_34_roi_V_reg  <= idata_34_roi_V;
      idata_35_roi_V_reg  <= idata_35_roi_V;
      idata_36_roi_V_reg  <= idata_36_roi_V;
      idata_37_roi_V_reg  <= idata_37_roi_V;
      idata_38_roi_V_reg  <= idata_38_roi_V;
      idata_39_roi_V_reg  <= idata_39_roi_V;
      idata_40_roi_V_reg  <= idata_40_roi_V;
      idata_41_roi_V_reg  <= idata_41_roi_V;
      idata_42_roi_V_reg  <= idata_42_roi_V;
      idata_43_roi_V_reg  <= idata_43_roi_V;
      idata_44_roi_V_reg  <= idata_44_roi_V;
      idata_45_roi_V_reg  <= idata_45_roi_V;
      idata_46_roi_V_reg  <= idata_46_roi_V;
      idata_47_roi_V_reg  <= idata_47_roi_V;
      idata_48_roi_V_reg  <= idata_48_roi_V;
      idata_49_roi_V_reg  <= idata_49_roi_V;
      idata_50_roi_V_reg  <= idata_50_roi_V;
      idata_51_roi_V_reg  <= idata_51_roi_V;
      idata_52_roi_V_reg  <= idata_52_roi_V;
      idata_53_roi_V_reg  <= idata_53_roi_V;
      idata_54_roi_V_reg  <= idata_54_roi_V;
      idata_55_roi_V_reg  <= idata_55_roi_V;
      idata_56_roi_V_reg  <= idata_56_roi_V;
      idata_57_roi_V_reg  <= idata_57_roi_V;
      idata_58_roi_V_reg  <= idata_58_roi_V;
      idata_59_roi_V_reg  <= idata_59_roi_V;
      idata_60_roi_V_reg  <= idata_60_roi_V;
      idata_61_roi_V_reg  <= idata_61_roi_V;
      idata_62_roi_V_reg  <= idata_62_roi_V;
      idata_63_roi_V_reg  <= idata_63_roi_V;
      idata_64_roi_V_reg  <= idata_64_roi_V;
      idata_65_roi_V_reg  <= idata_65_roi_V;
      idata_66_roi_V_reg  <= idata_66_roi_V;
      idata_67_roi_V_reg  <= idata_67_roi_V;
      idata_68_roi_V_reg  <= idata_68_roi_V;
      idata_69_roi_V_reg  <= idata_69_roi_V;
      idata_70_roi_V_reg  <= idata_70_roi_V;
      idata_71_roi_V_reg  <= idata_71_roi_V;
      idata_72_roi_V_reg  <= idata_72_roi_V;
      idata_73_roi_V_reg  <= idata_73_roi_V;
      idata_74_roi_V_reg  <= idata_74_roi_V;
      idata_75_roi_V_reg  <= idata_75_roi_V;
      idata_76_roi_V_reg  <= idata_76_roi_V;
      idata_77_roi_V_reg  <= idata_77_roi_V;
      idata_78_roi_V_reg  <= idata_78_roi_V;
      idata_79_roi_V_reg  <= idata_79_roi_V;
      idata_80_roi_V_reg  <= idata_80_roi_V;
      idata_81_roi_V_reg  <= idata_81_roi_V;
      idata_82_roi_V_reg  <= idata_82_roi_V;
      idata_83_roi_V_reg  <= idata_83_roi_V;
      idata_84_roi_V_reg  <= idata_84_roi_V;
      idata_85_roi_V_reg  <= idata_85_roi_V;
      idata_86_roi_V_reg  <= idata_86_roi_V;
      idata_87_roi_V_reg  <= idata_87_roi_V;
      idata_88_roi_V_reg  <= idata_88_roi_V;
      idata_89_roi_V_reg  <= idata_89_roi_V;
      idata_90_roi_V_reg  <= idata_90_roi_V;
      idata_91_roi_V_reg  <= idata_91_roi_V;
      idata_92_roi_V_reg  <= idata_92_roi_V;
      idata_93_roi_V_reg  <= idata_93_roi_V;
      idata_94_roi_V_reg  <= idata_94_roi_V;
      idata_95_roi_V_reg  <= idata_95_roi_V;
      idata_96_roi_V_reg  <= idata_96_roi_V;
      idata_97_roi_V_reg  <= idata_97_roi_V;
      idata_98_roi_V_reg  <= idata_98_roi_V;
      idata_99_roi_V_reg  <= idata_99_roi_V;
      idata_100_roi_V_reg <= idata_100_roi_V;
      idata_101_roi_V_reg <= idata_101_roi_V;
      idata_102_roi_V_reg <= idata_102_roi_V;
      idata_103_roi_V_reg <= idata_103_roi_V;
      idata_104_roi_V_reg <= idata_104_roi_V;
      idata_105_roi_V_reg <= idata_105_roi_V;
      idata_106_roi_V_reg <= idata_106_roi_V;
      idata_107_roi_V_reg <= idata_107_roi_V;
      idata_108_roi_V_reg <= idata_108_roi_V;
      idata_109_roi_V_reg <= idata_109_roi_V;
      idata_110_roi_V_reg <= idata_110_roi_V;
      idata_111_roi_V_reg <= idata_111_roi_V;
      idata_112_roi_V_reg <= idata_112_roi_V;
      idata_113_roi_V_reg <= idata_113_roi_V;
      idata_114_roi_V_reg <= idata_114_roi_V;
      idata_115_roi_V_reg <= idata_115_roi_V;
      idata_116_roi_V_reg <= idata_116_roi_V;
      idata_117_roi_V_reg <= idata_117_roi_V;
      idata_118_roi_V_reg <= idata_118_roi_V;
      idata_119_roi_V_reg <= idata_119_roi_V;
      idata_120_roi_V_reg <= idata_120_roi_V;
      idata_121_roi_V_reg <= idata_121_roi_V;
      idata_122_roi_V_reg <= idata_122_roi_V;
      idata_123_roi_V_reg <= idata_123_roi_V;
      idata_124_roi_V_reg <= idata_124_roi_V;
      idata_125_roi_V_reg <= idata_125_roi_V;
      idata_126_roi_V_reg <= idata_126_roi_V;
      idata_127_roi_V_reg <= idata_127_roi_V;
      idata_128_roi_V_reg <= idata_128_roi_V;
      idata_129_roi_V_reg <= idata_129_roi_V;
      idata_130_roi_V_reg <= idata_130_roi_V;
      idata_131_roi_V_reg <= idata_131_roi_V;
      idata_132_roi_V_reg <= idata_132_roi_V;
      idata_133_roi_V_reg <= idata_133_roi_V;
      idata_134_roi_V_reg <= idata_134_roi_V;
      idata_135_roi_V_reg <= idata_135_roi_V;
      idata_136_roi_V_reg <= idata_136_roi_V;
      idata_137_roi_V_reg <= idata_137_roi_V;
      idata_138_roi_V_reg <= idata_138_roi_V;
      idata_139_roi_V_reg <= idata_139_roi_V;
      idata_140_roi_V_reg <= idata_140_roi_V;
      idata_141_roi_V_reg <= idata_141_roi_V;
      idata_142_roi_V_reg <= idata_142_roi_V;
      idata_143_roi_V_reg <= idata_143_roi_V;
      idata_144_roi_V_reg <= idata_144_roi_V;
      idata_145_roi_V_reg <= idata_145_roi_V;
      idata_146_roi_V_reg <= idata_146_roi_V;
      idata_147_roi_V_reg <= idata_147_roi_V;
      idata_148_roi_V_reg <= idata_148_roi_V;
      idata_149_roi_V_reg <= idata_149_roi_V;
      idata_150_roi_V_reg <= idata_150_roi_V;
      idata_151_roi_V_reg <= idata_151_roi_V;
      idata_152_roi_V_reg <= idata_152_roi_V;
      idata_153_roi_V_reg <= idata_153_roi_V;
      idata_154_roi_V_reg <= idata_154_roi_V;
      idata_155_roi_V_reg <= idata_155_roi_V;
      idata_156_roi_V_reg <= idata_156_roi_V;
      idata_157_roi_V_reg <= idata_157_roi_V;
      idata_158_roi_V_reg <= idata_158_roi_V;
      idata_159_roi_V_reg <= idata_159_roi_V;
      idata_160_roi_V_reg <= idata_160_roi_V;
      idata_161_roi_V_reg <= idata_161_roi_V;
      idata_162_roi_V_reg <= idata_162_roi_V;
      idata_163_roi_V_reg <= idata_163_roi_V;
      idata_164_roi_V_reg <= idata_164_roi_V;
      idata_165_roi_V_reg <= idata_165_roi_V;
      idata_166_roi_V_reg <= idata_166_roi_V;
      idata_167_roi_V_reg <= idata_167_roi_V;
      idata_168_roi_V_reg <= idata_168_roi_V;
      idata_169_roi_V_reg <= idata_169_roi_V;
      idata_170_roi_V_reg <= idata_170_roi_V;
      idata_171_roi_V_reg <= idata_171_roi_V;
      idata_172_roi_V_reg <= idata_172_roi_V;
      idata_173_roi_V_reg <= idata_173_roi_V;
      idata_174_roi_V_reg <= idata_174_roi_V;
      idata_175_roi_V_reg <= idata_175_roi_V;
      idata_176_roi_V_reg <= idata_176_roi_V;
      idata_177_roi_V_reg <= idata_177_roi_V;
      idata_178_roi_V_reg <= idata_178_roi_V;
      idata_179_roi_V_reg <= idata_179_roi_V;
      idata_180_roi_V_reg <= idata_180_roi_V;
      idata_181_roi_V_reg <= idata_181_roi_V;
      idata_182_roi_V_reg <= idata_182_roi_V;
      idata_183_roi_V_reg <= idata_183_roi_V;
      idata_184_roi_V_reg <= idata_184_roi_V;
      idata_185_roi_V_reg <= idata_185_roi_V;
      idata_186_roi_V_reg <= idata_186_roi_V;
      idata_187_roi_V_reg <= idata_187_roi_V;
      idata_188_roi_V_reg <= idata_188_roi_V;
      idata_189_roi_V_reg <= idata_189_roi_V;
      idata_190_roi_V_reg <= idata_190_roi_V;
      idata_191_roi_V_reg <= idata_191_roi_V;
      idata_192_roi_V_reg <= idata_192_roi_V;
      idata_193_roi_V_reg <= idata_193_roi_V;
      idata_194_roi_V_reg <= idata_194_roi_V;
      idata_195_roi_V_reg <= idata_195_roi_V;
      idata_196_roi_V_reg <= idata_196_roi_V;
      idata_197_roi_V_reg <= idata_197_roi_V;
      idata_198_roi_V_reg <= idata_198_roi_V;
      idata_199_roi_V_reg <= idata_199_roi_V;
      idata_200_roi_V_reg <= idata_200_roi_V;
      idata_201_roi_V_reg <= idata_201_roi_V;
      idata_202_roi_V_reg <= idata_202_roi_V;
      idata_203_roi_V_reg <= idata_203_roi_V;
      idata_204_roi_V_reg <= idata_204_roi_V;
      idata_205_roi_V_reg <= idata_205_roi_V;
      idata_206_roi_V_reg <= idata_206_roi_V;
      idata_207_roi_V_reg <= idata_207_roi_V;
      idata_208_roi_V_reg <= idata_208_roi_V;
      idata_209_roi_V_reg <= idata_209_roi_V;
      idata_210_roi_V_reg <= idata_210_roi_V;
      idata_211_roi_V_reg <= idata_211_roi_V;
      idata_212_roi_V_reg <= idata_212_roi_V;
      idata_213_roi_V_reg <= idata_213_roi_V;
      idata_214_roi_V_reg <= idata_214_roi_V;
      idata_215_roi_V_reg <= idata_215_roi_V;
      idata_216_roi_V_reg <= idata_216_roi_V;
      idata_217_roi_V_reg <= idata_217_roi_V;
      idata_218_roi_V_reg <= idata_218_roi_V;
      idata_219_roi_V_reg <= idata_219_roi_V;
      idata_220_roi_V_reg <= idata_220_roi_V;
      idata_221_roi_V_reg <= idata_221_roi_V;
      idata_222_roi_V_reg <= idata_222_roi_V;
      idata_223_roi_V_reg <= idata_223_roi_V;
      idata_224_roi_V_reg <= idata_224_roi_V;
      idata_225_roi_V_reg <= idata_225_roi_V;
      idata_226_roi_V_reg <= idata_226_roi_V;
      idata_227_roi_V_reg <= idata_227_roi_V;
      idata_228_roi_V_reg <= idata_228_roi_V;
      idata_229_roi_V_reg <= idata_229_roi_V;
      idata_230_roi_V_reg <= idata_230_roi_V;
      idata_231_roi_V_reg <= idata_231_roi_V;
      idata_232_roi_V_reg <= idata_232_roi_V;
      idata_233_roi_V_reg <= idata_233_roi_V;
      idata_234_roi_V_reg <= idata_234_roi_V;
      idata_235_roi_V_reg <= idata_235_roi_V;
      idata_236_roi_V_reg <= idata_236_roi_V;
      idata_237_roi_V_reg <= idata_237_roi_V;
      idata_238_roi_V_reg <= idata_238_roi_V;
      idata_239_roi_V_reg <= idata_239_roi_V;
      idata_240_roi_V_reg <= idata_240_roi_V;
      idata_241_roi_V_reg <= idata_241_roi_V;
      idata_242_roi_V_reg <= idata_242_roi_V;
      idata_243_roi_V_reg <= idata_243_roi_V;
      idata_244_roi_V_reg <= idata_244_roi_V;
      idata_245_roi_V_reg <= idata_245_roi_V;
      idata_246_roi_V_reg <= idata_246_roi_V;
      idata_247_roi_V_reg <= idata_247_roi_V;
      idata_248_roi_V_reg <= idata_248_roi_V;
      idata_249_roi_V_reg <= idata_249_roi_V;
      idata_250_roi_V_reg <= idata_250_roi_V;
      idata_251_roi_V_reg <= idata_251_roi_V;
      idata_252_roi_V_reg <= idata_252_roi_V;
      idata_253_roi_V_reg <= idata_253_roi_V;
      idata_254_roi_V_reg <= idata_254_roi_V;
      idata_255_roi_V_reg <= idata_255_roi_V;
      idata_256_roi_V_reg <= idata_256_roi_V;
      idata_257_roi_V_reg <= idata_257_roi_V;
      idata_258_roi_V_reg <= idata_258_roi_V;
      idata_259_roi_V_reg <= idata_259_roi_V;
      idata_260_roi_V_reg <= idata_260_roi_V;
      idata_261_roi_V_reg <= idata_261_roi_V;
      idata_262_roi_V_reg <= idata_262_roi_V;
      idata_263_roi_V_reg <= idata_263_roi_V;
      idata_264_roi_V_reg <= idata_264_roi_V;
      idata_265_roi_V_reg <= idata_265_roi_V;
      idata_266_roi_V_reg <= idata_266_roi_V;
      idata_267_roi_V_reg <= idata_267_roi_V;
      idata_268_roi_V_reg <= idata_268_roi_V;
      idata_269_roi_V_reg <= idata_269_roi_V;
      idata_270_roi_V_reg <= idata_270_roi_V;
      idata_271_roi_V_reg <= idata_271_roi_V;
      idata_272_roi_V_reg <= idata_272_roi_V;
      idata_273_roi_V_reg <= idata_273_roi_V;
      idata_274_roi_V_reg <= idata_274_roi_V;
      idata_275_roi_V_reg <= idata_275_roi_V;
      idata_276_roi_V_reg <= idata_276_roi_V;
      idata_277_roi_V_reg <= idata_277_roi_V;
      idata_278_roi_V_reg <= idata_278_roi_V;
      idata_279_roi_V_reg <= idata_279_roi_V;
      idata_280_roi_V_reg <= idata_280_roi_V;
      idata_281_roi_V_reg <= idata_281_roi_V;
      idata_282_roi_V_reg <= idata_282_roi_V;
      idata_283_roi_V_reg <= idata_283_roi_V;
      idata_284_roi_V_reg <= idata_284_roi_V;
      idata_285_roi_V_reg <= idata_285_roi_V;
      idata_286_roi_V_reg <= idata_286_roi_V;
      idata_287_roi_V_reg <= idata_287_roi_V;
      idata_288_roi_V_reg <= idata_288_roi_V;
      idata_289_roi_V_reg <= idata_289_roi_V;
      idata_290_roi_V_reg <= idata_290_roi_V;
      idata_291_roi_V_reg <= idata_291_roi_V;
      idata_292_roi_V_reg <= idata_292_roi_V;
      idata_293_roi_V_reg <= idata_293_roi_V;
      idata_294_roi_V_reg <= idata_294_roi_V;
      idata_295_roi_V_reg <= idata_295_roi_V;
      idata_296_roi_V_reg <= idata_296_roi_V;
      idata_297_roi_V_reg <= idata_297_roi_V;
      idata_298_roi_V_reg <= idata_298_roi_V;
      idata_299_roi_V_reg <= idata_299_roi_V;
      idata_300_roi_V_reg <= idata_300_roi_V;
      idata_301_roi_V_reg <= idata_301_roi_V;
      idata_302_roi_V_reg <= idata_302_roi_V;
      idata_303_roi_V_reg <= idata_303_roi_V;
      idata_304_roi_V_reg <= idata_304_roi_V;
      idata_305_roi_V_reg <= idata_305_roi_V;
      idata_306_roi_V_reg <= idata_306_roi_V;
      idata_307_roi_V_reg <= idata_307_roi_V;
      idata_308_roi_V_reg <= idata_308_roi_V;
      idata_309_roi_V_reg <= idata_309_roi_V;
      idata_310_roi_V_reg <= idata_310_roi_V;
      idata_311_roi_V_reg <= idata_311_roi_V;
      idata_312_roi_V_reg <= idata_312_roi_V;
      idata_313_roi_V_reg <= idata_313_roi_V;
      idata_314_roi_V_reg <= idata_314_roi_V;
      idata_315_roi_V_reg <= idata_315_roi_V;
      idata_316_roi_V_reg <= idata_316_roi_V;
      idata_317_roi_V_reg <= idata_317_roi_V;
      idata_318_roi_V_reg <= idata_318_roi_V;
      idata_319_roi_V_reg <= idata_319_roi_V;
      idata_320_roi_V_reg <= idata_320_roi_V;
      idata_321_roi_V_reg <= idata_321_roi_V;
      idata_322_roi_V_reg <= idata_322_roi_V;
      idata_323_roi_V_reg <= idata_323_roi_V;
      idata_324_roi_V_reg <= idata_324_roi_V;
      idata_325_roi_V_reg <= idata_325_roi_V;
      idata_326_roi_V_reg <= idata_326_roi_V;
      idata_327_roi_V_reg <= idata_327_roi_V;
      idata_328_roi_V_reg <= idata_328_roi_V;
      idata_329_roi_V_reg <= idata_329_roi_V;
      idata_330_roi_V_reg <= idata_330_roi_V;
      idata_331_roi_V_reg <= idata_331_roi_V;
      idata_332_roi_V_reg <= idata_332_roi_V;
      idata_333_roi_V_reg <= idata_333_roi_V;
      idata_334_roi_V_reg <= idata_334_roi_V;
      idata_335_roi_V_reg <= idata_335_roi_V;
      idata_336_roi_V_reg <= idata_336_roi_V;
      idata_337_roi_V_reg <= idata_337_roi_V;
      idata_338_roi_V_reg <= idata_338_roi_V;
      idata_339_roi_V_reg <= idata_339_roi_V;
      idata_340_roi_V_reg <= idata_340_roi_V;
      idata_341_roi_V_reg <= idata_341_roi_V;
      idata_342_roi_V_reg <= idata_342_roi_V;
      idata_343_roi_V_reg <= idata_343_roi_V;
      idata_344_roi_V_reg <= idata_344_roi_V;
      idata_345_roi_V_reg <= idata_345_roi_V;
      idata_346_roi_V_reg <= idata_346_roi_V;
      idata_347_roi_V_reg <= idata_347_roi_V;
      idata_348_roi_V_reg <= idata_348_roi_V;
      idata_349_roi_V_reg <= idata_349_roi_V;
      idata_350_roi_V_reg <= idata_350_roi_V;
      idata_351_roi_V_reg <= idata_351_roi_V;
      idata_0_flg_V_reg   <= idata_0_flg_V;
      idata_1_flg_V_reg   <= idata_1_flg_V;
      idata_2_flg_V_reg   <= idata_2_flg_V;
      idata_3_flg_V_reg   <= idata_3_flg_V;
      idata_4_flg_V_reg   <= idata_4_flg_V;
      idata_5_flg_V_reg   <= idata_5_flg_V;
      idata_6_flg_V_reg   <= idata_6_flg_V;
      idata_7_flg_V_reg   <= idata_7_flg_V;
      idata_8_flg_V_reg   <= idata_8_flg_V;
      idata_9_flg_V_reg   <= idata_9_flg_V;
      idata_10_flg_V_reg  <= idata_10_flg_V;
      idata_11_flg_V_reg  <= idata_11_flg_V;
      idata_12_flg_V_reg  <= idata_12_flg_V;
      idata_13_flg_V_reg  <= idata_13_flg_V;
      idata_14_flg_V_reg  <= idata_14_flg_V;
      idata_15_flg_V_reg  <= idata_15_flg_V;
      idata_16_flg_V_reg  <= idata_16_flg_V;
      idata_17_flg_V_reg  <= idata_17_flg_V;
      idata_18_flg_V_reg  <= idata_18_flg_V;
      idata_19_flg_V_reg  <= idata_19_flg_V;
      idata_20_flg_V_reg  <= idata_20_flg_V;
      idata_21_flg_V_reg  <= idata_21_flg_V;
      idata_22_flg_V_reg  <= idata_22_flg_V;
      idata_23_flg_V_reg  <= idata_23_flg_V;
      idata_24_flg_V_reg  <= idata_24_flg_V;
      idata_25_flg_V_reg  <= idata_25_flg_V;
      idata_26_flg_V_reg  <= idata_26_flg_V;
      idata_27_flg_V_reg  <= idata_27_flg_V;
      idata_28_flg_V_reg  <= idata_28_flg_V;
      idata_29_flg_V_reg  <= idata_29_flg_V;
      idata_30_flg_V_reg  <= idata_30_flg_V;
      idata_31_flg_V_reg  <= idata_31_flg_V;
      idata_32_flg_V_reg  <= idata_32_flg_V;
      idata_33_flg_V_reg  <= idata_33_flg_V;
      idata_34_flg_V_reg  <= idata_34_flg_V;
      idata_35_flg_V_reg  <= idata_35_flg_V;
      idata_36_flg_V_reg  <= idata_36_flg_V;
      idata_37_flg_V_reg  <= idata_37_flg_V;
      idata_38_flg_V_reg  <= idata_38_flg_V;
      idata_39_flg_V_reg  <= idata_39_flg_V;
      idata_40_flg_V_reg  <= idata_40_flg_V;
      idata_41_flg_V_reg  <= idata_41_flg_V;
      idata_42_flg_V_reg  <= idata_42_flg_V;
      idata_43_flg_V_reg  <= idata_43_flg_V;
      idata_44_flg_V_reg  <= idata_44_flg_V;
      idata_45_flg_V_reg  <= idata_45_flg_V;
      idata_46_flg_V_reg  <= idata_46_flg_V;
      idata_47_flg_V_reg  <= idata_47_flg_V;
      idata_48_flg_V_reg  <= idata_48_flg_V;
      idata_49_flg_V_reg  <= idata_49_flg_V;
      idata_50_flg_V_reg  <= idata_50_flg_V;
      idata_51_flg_V_reg  <= idata_51_flg_V;
      idata_52_flg_V_reg  <= idata_52_flg_V;
      idata_53_flg_V_reg  <= idata_53_flg_V;
      idata_54_flg_V_reg  <= idata_54_flg_V;
      idata_55_flg_V_reg  <= idata_55_flg_V;
      idata_56_flg_V_reg  <= idata_56_flg_V;
      idata_57_flg_V_reg  <= idata_57_flg_V;
      idata_58_flg_V_reg  <= idata_58_flg_V;
      idata_59_flg_V_reg  <= idata_59_flg_V;
      idata_60_flg_V_reg  <= idata_60_flg_V;
      idata_61_flg_V_reg  <= idata_61_flg_V;
      idata_62_flg_V_reg  <= idata_62_flg_V;
      idata_63_flg_V_reg  <= idata_63_flg_V;
      idata_64_flg_V_reg  <= idata_64_flg_V;
      idata_65_flg_V_reg  <= idata_65_flg_V;
      idata_66_flg_V_reg  <= idata_66_flg_V;
      idata_67_flg_V_reg  <= idata_67_flg_V;
      idata_68_flg_V_reg  <= idata_68_flg_V;
      idata_69_flg_V_reg  <= idata_69_flg_V;
      idata_70_flg_V_reg  <= idata_70_flg_V;
      idata_71_flg_V_reg  <= idata_71_flg_V;
      idata_72_flg_V_reg  <= idata_72_flg_V;
      idata_73_flg_V_reg  <= idata_73_flg_V;
      idata_74_flg_V_reg  <= idata_74_flg_V;
      idata_75_flg_V_reg  <= idata_75_flg_V;
      idata_76_flg_V_reg  <= idata_76_flg_V;
      idata_77_flg_V_reg  <= idata_77_flg_V;
      idata_78_flg_V_reg  <= idata_78_flg_V;
      idata_79_flg_V_reg  <= idata_79_flg_V;
      idata_80_flg_V_reg  <= idata_80_flg_V;
      idata_81_flg_V_reg  <= idata_81_flg_V;
      idata_82_flg_V_reg  <= idata_82_flg_V;
      idata_83_flg_V_reg  <= idata_83_flg_V;
      idata_84_flg_V_reg  <= idata_84_flg_V;
      idata_85_flg_V_reg  <= idata_85_flg_V;
      idata_86_flg_V_reg  <= idata_86_flg_V;
      idata_87_flg_V_reg  <= idata_87_flg_V;
      idata_88_flg_V_reg  <= idata_88_flg_V;
      idata_89_flg_V_reg  <= idata_89_flg_V;
      idata_90_flg_V_reg  <= idata_90_flg_V;
      idata_91_flg_V_reg  <= idata_91_flg_V;
      idata_92_flg_V_reg  <= idata_92_flg_V;
      idata_93_flg_V_reg  <= idata_93_flg_V;
      idata_94_flg_V_reg  <= idata_94_flg_V;
      idata_95_flg_V_reg  <= idata_95_flg_V;
      idata_96_flg_V_reg  <= idata_96_flg_V;
      idata_97_flg_V_reg  <= idata_97_flg_V;
      idata_98_flg_V_reg  <= idata_98_flg_V;
      idata_99_flg_V_reg  <= idata_99_flg_V;
      idata_100_flg_V_reg <= idata_100_flg_V;
      idata_101_flg_V_reg <= idata_101_flg_V;
      idata_102_flg_V_reg <= idata_102_flg_V;
      idata_103_flg_V_reg <= idata_103_flg_V;
      idata_104_flg_V_reg <= idata_104_flg_V;
      idata_105_flg_V_reg <= idata_105_flg_V;
      idata_106_flg_V_reg <= idata_106_flg_V;
      idata_107_flg_V_reg <= idata_107_flg_V;
      idata_108_flg_V_reg <= idata_108_flg_V;
      idata_109_flg_V_reg <= idata_109_flg_V;
      idata_110_flg_V_reg <= idata_110_flg_V;
      idata_111_flg_V_reg <= idata_111_flg_V;
      idata_112_flg_V_reg <= idata_112_flg_V;
      idata_113_flg_V_reg <= idata_113_flg_V;
      idata_114_flg_V_reg <= idata_114_flg_V;
      idata_115_flg_V_reg <= idata_115_flg_V;
      idata_116_flg_V_reg <= idata_116_flg_V;
      idata_117_flg_V_reg <= idata_117_flg_V;
      idata_118_flg_V_reg <= idata_118_flg_V;
      idata_119_flg_V_reg <= idata_119_flg_V;
      idata_120_flg_V_reg <= idata_120_flg_V;
      idata_121_flg_V_reg <= idata_121_flg_V;
      idata_122_flg_V_reg <= idata_122_flg_V;
      idata_123_flg_V_reg <= idata_123_flg_V;
      idata_124_flg_V_reg <= idata_124_flg_V;
      idata_125_flg_V_reg <= idata_125_flg_V;
      idata_126_flg_V_reg <= idata_126_flg_V;
      idata_127_flg_V_reg <= idata_127_flg_V;
      idata_128_flg_V_reg <= idata_128_flg_V;
      idata_129_flg_V_reg <= idata_129_flg_V;
      idata_130_flg_V_reg <= idata_130_flg_V;
      idata_131_flg_V_reg <= idata_131_flg_V;
      idata_132_flg_V_reg <= idata_132_flg_V;
      idata_133_flg_V_reg <= idata_133_flg_V;
      idata_134_flg_V_reg <= idata_134_flg_V;
      idata_135_flg_V_reg <= idata_135_flg_V;
      idata_136_flg_V_reg <= idata_136_flg_V;
      idata_137_flg_V_reg <= idata_137_flg_V;
      idata_138_flg_V_reg <= idata_138_flg_V;
      idata_139_flg_V_reg <= idata_139_flg_V;
      idata_140_flg_V_reg <= idata_140_flg_V;
      idata_141_flg_V_reg <= idata_141_flg_V;
      idata_142_flg_V_reg <= idata_142_flg_V;
      idata_143_flg_V_reg <= idata_143_flg_V;
      idata_144_flg_V_reg <= idata_144_flg_V;
      idata_145_flg_V_reg <= idata_145_flg_V;
      idata_146_flg_V_reg <= idata_146_flg_V;
      idata_147_flg_V_reg <= idata_147_flg_V;
      idata_148_flg_V_reg <= idata_148_flg_V;
      idata_149_flg_V_reg <= idata_149_flg_V;
      idata_150_flg_V_reg <= idata_150_flg_V;
      idata_151_flg_V_reg <= idata_151_flg_V;
      idata_152_flg_V_reg <= idata_152_flg_V;
      idata_153_flg_V_reg <= idata_153_flg_V;
      idata_154_flg_V_reg <= idata_154_flg_V;
      idata_155_flg_V_reg <= idata_155_flg_V;
      idata_156_flg_V_reg <= idata_156_flg_V;
      idata_157_flg_V_reg <= idata_157_flg_V;
      idata_158_flg_V_reg <= idata_158_flg_V;
      idata_159_flg_V_reg <= idata_159_flg_V;
      idata_160_flg_V_reg <= idata_160_flg_V;
      idata_161_flg_V_reg <= idata_161_flg_V;
      idata_162_flg_V_reg <= idata_162_flg_V;
      idata_163_flg_V_reg <= idata_163_flg_V;
      idata_164_flg_V_reg <= idata_164_flg_V;
      idata_165_flg_V_reg <= idata_165_flg_V;
      idata_166_flg_V_reg <= idata_166_flg_V;
      idata_167_flg_V_reg <= idata_167_flg_V;
      idata_168_flg_V_reg <= idata_168_flg_V;
      idata_169_flg_V_reg <= idata_169_flg_V;
      idata_170_flg_V_reg <= idata_170_flg_V;
      idata_171_flg_V_reg <= idata_171_flg_V;
      idata_172_flg_V_reg <= idata_172_flg_V;
      idata_173_flg_V_reg <= idata_173_flg_V;
      idata_174_flg_V_reg <= idata_174_flg_V;
      idata_175_flg_V_reg <= idata_175_flg_V;
      idata_176_flg_V_reg <= idata_176_flg_V;
      idata_177_flg_V_reg <= idata_177_flg_V;
      idata_178_flg_V_reg <= idata_178_flg_V;
      idata_179_flg_V_reg <= idata_179_flg_V;
      idata_180_flg_V_reg <= idata_180_flg_V;
      idata_181_flg_V_reg <= idata_181_flg_V;
      idata_182_flg_V_reg <= idata_182_flg_V;
      idata_183_flg_V_reg <= idata_183_flg_V;
      idata_184_flg_V_reg <= idata_184_flg_V;
      idata_185_flg_V_reg <= idata_185_flg_V;
      idata_186_flg_V_reg <= idata_186_flg_V;
      idata_187_flg_V_reg <= idata_187_flg_V;
      idata_188_flg_V_reg <= idata_188_flg_V;
      idata_189_flg_V_reg <= idata_189_flg_V;
      idata_190_flg_V_reg <= idata_190_flg_V;
      idata_191_flg_V_reg <= idata_191_flg_V;
      idata_192_flg_V_reg <= idata_192_flg_V;
      idata_193_flg_V_reg <= idata_193_flg_V;
      idata_194_flg_V_reg <= idata_194_flg_V;
      idata_195_flg_V_reg <= idata_195_flg_V;
      idata_196_flg_V_reg <= idata_196_flg_V;
      idata_197_flg_V_reg <= idata_197_flg_V;
      idata_198_flg_V_reg <= idata_198_flg_V;
      idata_199_flg_V_reg <= idata_199_flg_V;
      idata_200_flg_V_reg <= idata_200_flg_V;
      idata_201_flg_V_reg <= idata_201_flg_V;
      idata_202_flg_V_reg <= idata_202_flg_V;
      idata_203_flg_V_reg <= idata_203_flg_V;
      idata_204_flg_V_reg <= idata_204_flg_V;
      idata_205_flg_V_reg <= idata_205_flg_V;
      idata_206_flg_V_reg <= idata_206_flg_V;
      idata_207_flg_V_reg <= idata_207_flg_V;
      idata_208_flg_V_reg <= idata_208_flg_V;
      idata_209_flg_V_reg <= idata_209_flg_V;
      idata_210_flg_V_reg <= idata_210_flg_V;
      idata_211_flg_V_reg <= idata_211_flg_V;
      idata_212_flg_V_reg <= idata_212_flg_V;
      idata_213_flg_V_reg <= idata_213_flg_V;
      idata_214_flg_V_reg <= idata_214_flg_V;
      idata_215_flg_V_reg <= idata_215_flg_V;
      idata_216_flg_V_reg <= idata_216_flg_V;
      idata_217_flg_V_reg <= idata_217_flg_V;
      idata_218_flg_V_reg <= idata_218_flg_V;
      idata_219_flg_V_reg <= idata_219_flg_V;
      idata_220_flg_V_reg <= idata_220_flg_V;
      idata_221_flg_V_reg <= idata_221_flg_V;
      idata_222_flg_V_reg <= idata_222_flg_V;
      idata_223_flg_V_reg <= idata_223_flg_V;
      idata_224_flg_V_reg <= idata_224_flg_V;
      idata_225_flg_V_reg <= idata_225_flg_V;
      idata_226_flg_V_reg <= idata_226_flg_V;
      idata_227_flg_V_reg <= idata_227_flg_V;
      idata_228_flg_V_reg <= idata_228_flg_V;
      idata_229_flg_V_reg <= idata_229_flg_V;
      idata_230_flg_V_reg <= idata_230_flg_V;
      idata_231_flg_V_reg <= idata_231_flg_V;
      idata_232_flg_V_reg <= idata_232_flg_V;
      idata_233_flg_V_reg <= idata_233_flg_V;
      idata_234_flg_V_reg <= idata_234_flg_V;
      idata_235_flg_V_reg <= idata_235_flg_V;
      idata_236_flg_V_reg <= idata_236_flg_V;
      idata_237_flg_V_reg <= idata_237_flg_V;
      idata_238_flg_V_reg <= idata_238_flg_V;
      idata_239_flg_V_reg <= idata_239_flg_V;
      idata_240_flg_V_reg <= idata_240_flg_V;
      idata_241_flg_V_reg <= idata_241_flg_V;
      idata_242_flg_V_reg <= idata_242_flg_V;
      idata_243_flg_V_reg <= idata_243_flg_V;
      idata_244_flg_V_reg <= idata_244_flg_V;
      idata_245_flg_V_reg <= idata_245_flg_V;
      idata_246_flg_V_reg <= idata_246_flg_V;
      idata_247_flg_V_reg <= idata_247_flg_V;
      idata_248_flg_V_reg <= idata_248_flg_V;
      idata_249_flg_V_reg <= idata_249_flg_V;
      idata_250_flg_V_reg <= idata_250_flg_V;
      idata_251_flg_V_reg <= idata_251_flg_V;
      idata_252_flg_V_reg <= idata_252_flg_V;
      idata_253_flg_V_reg <= idata_253_flg_V;
      idata_254_flg_V_reg <= idata_254_flg_V;
      idata_255_flg_V_reg <= idata_255_flg_V;
      idata_256_flg_V_reg <= idata_256_flg_V;
      idata_257_flg_V_reg <= idata_257_flg_V;
      idata_258_flg_V_reg <= idata_258_flg_V;
      idata_259_flg_V_reg <= idata_259_flg_V;
      idata_260_flg_V_reg <= idata_260_flg_V;
      idata_261_flg_V_reg <= idata_261_flg_V;
      idata_262_flg_V_reg <= idata_262_flg_V;
      idata_263_flg_V_reg <= idata_263_flg_V;
      idata_264_flg_V_reg <= idata_264_flg_V;
      idata_265_flg_V_reg <= idata_265_flg_V;
      idata_266_flg_V_reg <= idata_266_flg_V;
      idata_267_flg_V_reg <= idata_267_flg_V;
      idata_268_flg_V_reg <= idata_268_flg_V;
      idata_269_flg_V_reg <= idata_269_flg_V;
      idata_270_flg_V_reg <= idata_270_flg_V;
      idata_271_flg_V_reg <= idata_271_flg_V;
      idata_272_flg_V_reg <= idata_272_flg_V;
      idata_273_flg_V_reg <= idata_273_flg_V;
      idata_274_flg_V_reg <= idata_274_flg_V;
      idata_275_flg_V_reg <= idata_275_flg_V;
      idata_276_flg_V_reg <= idata_276_flg_V;
      idata_277_flg_V_reg <= idata_277_flg_V;
      idata_278_flg_V_reg <= idata_278_flg_V;
      idata_279_flg_V_reg <= idata_279_flg_V;
      idata_280_flg_V_reg <= idata_280_flg_V;
      idata_281_flg_V_reg <= idata_281_flg_V;
      idata_282_flg_V_reg <= idata_282_flg_V;
      idata_283_flg_V_reg <= idata_283_flg_V;
      idata_284_flg_V_reg <= idata_284_flg_V;
      idata_285_flg_V_reg <= idata_285_flg_V;
      idata_286_flg_V_reg <= idata_286_flg_V;
      idata_287_flg_V_reg <= idata_287_flg_V;
      idata_288_flg_V_reg <= idata_288_flg_V;
      idata_289_flg_V_reg <= idata_289_flg_V;
      idata_290_flg_V_reg <= idata_290_flg_V;
      idata_291_flg_V_reg <= idata_291_flg_V;
      idata_292_flg_V_reg <= idata_292_flg_V;
      idata_293_flg_V_reg <= idata_293_flg_V;
      idata_294_flg_V_reg <= idata_294_flg_V;
      idata_295_flg_V_reg <= idata_295_flg_V;
      idata_296_flg_V_reg <= idata_296_flg_V;
      idata_297_flg_V_reg <= idata_297_flg_V;
      idata_298_flg_V_reg <= idata_298_flg_V;
      idata_299_flg_V_reg <= idata_299_flg_V;
      idata_300_flg_V_reg <= idata_300_flg_V;
      idata_301_flg_V_reg <= idata_301_flg_V;
      idata_302_flg_V_reg <= idata_302_flg_V;
      idata_303_flg_V_reg <= idata_303_flg_V;
      idata_304_flg_V_reg <= idata_304_flg_V;
      idata_305_flg_V_reg <= idata_305_flg_V;
      idata_306_flg_V_reg <= idata_306_flg_V;
      idata_307_flg_V_reg <= idata_307_flg_V;
      idata_308_flg_V_reg <= idata_308_flg_V;
      idata_309_flg_V_reg <= idata_309_flg_V;
      idata_310_flg_V_reg <= idata_310_flg_V;
      idata_311_flg_V_reg <= idata_311_flg_V;
      idata_312_flg_V_reg <= idata_312_flg_V;
      idata_313_flg_V_reg <= idata_313_flg_V;
      idata_314_flg_V_reg <= idata_314_flg_V;
      idata_315_flg_V_reg <= idata_315_flg_V;
      idata_316_flg_V_reg <= idata_316_flg_V;
      idata_317_flg_V_reg <= idata_317_flg_V;
      idata_318_flg_V_reg <= idata_318_flg_V;
      idata_319_flg_V_reg <= idata_319_flg_V;
      idata_320_flg_V_reg <= idata_320_flg_V;
      idata_321_flg_V_reg <= idata_321_flg_V;
      idata_322_flg_V_reg <= idata_322_flg_V;
      idata_323_flg_V_reg <= idata_323_flg_V;
      idata_324_flg_V_reg <= idata_324_flg_V;
      idata_325_flg_V_reg <= idata_325_flg_V;
      idata_326_flg_V_reg <= idata_326_flg_V;
      idata_327_flg_V_reg <= idata_327_flg_V;
      idata_328_flg_V_reg <= idata_328_flg_V;
      idata_329_flg_V_reg <= idata_329_flg_V;
      idata_330_flg_V_reg <= idata_330_flg_V;
      idata_331_flg_V_reg <= idata_331_flg_V;
      idata_332_flg_V_reg <= idata_332_flg_V;
      idata_333_flg_V_reg <= idata_333_flg_V;
      idata_334_flg_V_reg <= idata_334_flg_V;
      idata_335_flg_V_reg <= idata_335_flg_V;
      idata_336_flg_V_reg <= idata_336_flg_V;
      idata_337_flg_V_reg <= idata_337_flg_V;
      idata_338_flg_V_reg <= idata_338_flg_V;
      idata_339_flg_V_reg <= idata_339_flg_V;
      idata_340_flg_V_reg <= idata_340_flg_V;
      idata_341_flg_V_reg <= idata_341_flg_V;
      idata_342_flg_V_reg <= idata_342_flg_V;
      idata_343_flg_V_reg <= idata_343_flg_V;
      idata_344_flg_V_reg <= idata_344_flg_V;
      idata_345_flg_V_reg <= idata_345_flg_V;
      idata_346_flg_V_reg <= idata_346_flg_V;
      idata_347_flg_V_reg <= idata_347_flg_V;
      idata_348_flg_V_reg <= idata_348_flg_V;
      idata_349_flg_V_reg <= idata_349_flg_V;
      idata_350_flg_V_reg <= idata_350_flg_V;
      idata_351_flg_V_reg <= idata_351_flg_V;

      
    end if;
  end process reg_p;




  -- DUT

  compare_main_1 : component compare_main
    port map (
      ap_clk          => ap_clk,
      ap_rst          => ap_rst,
      ap_start        => ap_start_reg,
      ap_done         => ap_done,
      ap_idle         => ap_idle,
      ap_ready        => ap_ready,
      idata_0_pt_V    => idata_0_pt_V_reg,
      idata_1_pt_V    => idata_1_pt_V_reg,
      idata_2_pt_V    => idata_2_pt_V_reg,
      idata_3_pt_V    => idata_3_pt_V_reg,
      idata_4_pt_V    => idata_4_pt_V_reg,
      idata_5_pt_V    => idata_5_pt_V_reg,
      idata_6_pt_V    => idata_6_pt_V_reg,
      idata_7_pt_V    => idata_7_pt_V_reg,
      idata_8_pt_V    => idata_8_pt_V_reg,
      idata_9_pt_V    => idata_9_pt_V_reg,
      idata_10_pt_V   => idata_10_pt_V_reg,
      idata_11_pt_V   => idata_11_pt_V_reg,
      idata_12_pt_V   => idata_12_pt_V_reg,
      idata_13_pt_V   => idata_13_pt_V_reg,
      idata_14_pt_V   => idata_14_pt_V_reg,
      idata_15_pt_V   => idata_15_pt_V_reg,
      idata_16_pt_V   => idata_16_pt_V_reg,
      idata_17_pt_V   => idata_17_pt_V_reg,
      idata_18_pt_V   => idata_18_pt_V_reg,
      idata_19_pt_V   => idata_19_pt_V_reg,
      idata_20_pt_V   => idata_20_pt_V_reg,
      idata_21_pt_V   => idata_21_pt_V_reg,
      idata_22_pt_V   => idata_22_pt_V_reg,
      idata_23_pt_V   => idata_23_pt_V_reg,
      idata_24_pt_V   => idata_24_pt_V_reg,
      idata_25_pt_V   => idata_25_pt_V_reg,
      idata_26_pt_V   => idata_26_pt_V_reg,
      idata_27_pt_V   => idata_27_pt_V_reg,
      idata_28_pt_V   => idata_28_pt_V_reg,
      idata_29_pt_V   => idata_29_pt_V_reg,
      idata_30_pt_V   => idata_30_pt_V_reg,
      idata_31_pt_V   => idata_31_pt_V_reg,
      idata_32_pt_V   => idata_32_pt_V_reg,
      idata_33_pt_V   => idata_33_pt_V_reg,
      idata_34_pt_V   => idata_34_pt_V_reg,
      idata_35_pt_V   => idata_35_pt_V_reg,
      idata_36_pt_V   => idata_36_pt_V_reg,
      idata_37_pt_V   => idata_37_pt_V_reg,
      idata_38_pt_V   => idata_38_pt_V_reg,
      idata_39_pt_V   => idata_39_pt_V_reg,
      idata_40_pt_V   => idata_40_pt_V_reg,
      idata_41_pt_V   => idata_41_pt_V_reg,
      idata_42_pt_V   => idata_42_pt_V_reg,
      idata_43_pt_V   => idata_43_pt_V_reg,
      idata_44_pt_V   => idata_44_pt_V_reg,
      idata_45_pt_V   => idata_45_pt_V_reg,
      idata_46_pt_V   => idata_46_pt_V_reg,
      idata_47_pt_V   => idata_47_pt_V_reg,
      idata_48_pt_V   => idata_48_pt_V_reg,
      idata_49_pt_V   => idata_49_pt_V_reg,
      idata_50_pt_V   => idata_50_pt_V_reg,
      idata_51_pt_V   => idata_51_pt_V_reg,
      idata_52_pt_V   => idata_52_pt_V_reg,
      idata_53_pt_V   => idata_53_pt_V_reg,
      idata_54_pt_V   => idata_54_pt_V_reg,
      idata_55_pt_V   => idata_55_pt_V_reg,
      idata_56_pt_V   => idata_56_pt_V_reg,
      idata_57_pt_V   => idata_57_pt_V_reg,
      idata_58_pt_V   => idata_58_pt_V_reg,
      idata_59_pt_V   => idata_59_pt_V_reg,
      idata_60_pt_V   => idata_60_pt_V_reg,
      idata_61_pt_V   => idata_61_pt_V_reg,
      idata_62_pt_V   => idata_62_pt_V_reg,
      idata_63_pt_V   => idata_63_pt_V_reg,
      idata_64_pt_V   => idata_64_pt_V_reg,
      idata_65_pt_V   => idata_65_pt_V_reg,
      idata_66_pt_V   => idata_66_pt_V_reg,
      idata_67_pt_V   => idata_67_pt_V_reg,
      idata_68_pt_V   => idata_68_pt_V_reg,
      idata_69_pt_V   => idata_69_pt_V_reg,
      idata_70_pt_V   => idata_70_pt_V_reg,
      idata_71_pt_V   => idata_71_pt_V_reg,
      idata_72_pt_V   => idata_72_pt_V_reg,
      idata_73_pt_V   => idata_73_pt_V_reg,
      idata_74_pt_V   => idata_74_pt_V_reg,
      idata_75_pt_V   => idata_75_pt_V_reg,
      idata_76_pt_V   => idata_76_pt_V_reg,
      idata_77_pt_V   => idata_77_pt_V_reg,
      idata_78_pt_V   => idata_78_pt_V_reg,
      idata_79_pt_V   => idata_79_pt_V_reg,
      idata_80_pt_V   => idata_80_pt_V_reg,
      idata_81_pt_V   => idata_81_pt_V_reg,
      idata_82_pt_V   => idata_82_pt_V_reg,
      idata_83_pt_V   => idata_83_pt_V_reg,
      idata_84_pt_V   => idata_84_pt_V_reg,
      idata_85_pt_V   => idata_85_pt_V_reg,
      idata_86_pt_V   => idata_86_pt_V_reg,
      idata_87_pt_V   => idata_87_pt_V_reg,
      idata_88_pt_V   => idata_88_pt_V_reg,
      idata_89_pt_V   => idata_89_pt_V_reg,
      idata_90_pt_V   => idata_90_pt_V_reg,
      idata_91_pt_V   => idata_91_pt_V_reg,
      idata_92_pt_V   => idata_92_pt_V_reg,
      idata_93_pt_V   => idata_93_pt_V_reg,
      idata_94_pt_V   => idata_94_pt_V_reg,
      idata_95_pt_V   => idata_95_pt_V_reg,
      idata_96_pt_V   => idata_96_pt_V_reg,
      idata_97_pt_V   => idata_97_pt_V_reg,
      idata_98_pt_V   => idata_98_pt_V_reg,
      idata_99_pt_V   => idata_99_pt_V_reg,
      idata_100_pt_V  => idata_100_pt_V_reg,
      idata_101_pt_V  => idata_101_pt_V_reg,
      idata_102_pt_V  => idata_102_pt_V_reg,
      idata_103_pt_V  => idata_103_pt_V_reg,
      idata_104_pt_V  => idata_104_pt_V_reg,
      idata_105_pt_V  => idata_105_pt_V_reg,
      idata_106_pt_V  => idata_106_pt_V_reg,
      idata_107_pt_V  => idata_107_pt_V_reg,
      idata_108_pt_V  => idata_108_pt_V_reg,
      idata_109_pt_V  => idata_109_pt_V_reg,
      idata_110_pt_V  => idata_110_pt_V_reg,
      idata_111_pt_V  => idata_111_pt_V_reg,
      idata_112_pt_V  => idata_112_pt_V_reg,
      idata_113_pt_V  => idata_113_pt_V_reg,
      idata_114_pt_V  => idata_114_pt_V_reg,
      idata_115_pt_V  => idata_115_pt_V_reg,
      idata_116_pt_V  => idata_116_pt_V_reg,
      idata_117_pt_V  => idata_117_pt_V_reg,
      idata_118_pt_V  => idata_118_pt_V_reg,
      idata_119_pt_V  => idata_119_pt_V_reg,
      idata_120_pt_V  => idata_120_pt_V_reg,
      idata_121_pt_V  => idata_121_pt_V_reg,
      idata_122_pt_V  => idata_122_pt_V_reg,
      idata_123_pt_V  => idata_123_pt_V_reg,
      idata_124_pt_V  => idata_124_pt_V_reg,
      idata_125_pt_V  => idata_125_pt_V_reg,
      idata_126_pt_V  => idata_126_pt_V_reg,
      idata_127_pt_V  => idata_127_pt_V_reg,
      idata_128_pt_V  => idata_128_pt_V_reg,
      idata_129_pt_V  => idata_129_pt_V_reg,
      idata_130_pt_V  => idata_130_pt_V_reg,
      idata_131_pt_V  => idata_131_pt_V_reg,
      idata_132_pt_V  => idata_132_pt_V_reg,
      idata_133_pt_V  => idata_133_pt_V_reg,
      idata_134_pt_V  => idata_134_pt_V_reg,
      idata_135_pt_V  => idata_135_pt_V_reg,
      idata_136_pt_V  => idata_136_pt_V_reg,
      idata_137_pt_V  => idata_137_pt_V_reg,
      idata_138_pt_V  => idata_138_pt_V_reg,
      idata_139_pt_V  => idata_139_pt_V_reg,
      idata_140_pt_V  => idata_140_pt_V_reg,
      idata_141_pt_V  => idata_141_pt_V_reg,
      idata_142_pt_V  => idata_142_pt_V_reg,
      idata_143_pt_V  => idata_143_pt_V_reg,
      idata_144_pt_V  => idata_144_pt_V_reg,
      idata_145_pt_V  => idata_145_pt_V_reg,
      idata_146_pt_V  => idata_146_pt_V_reg,
      idata_147_pt_V  => idata_147_pt_V_reg,
      idata_148_pt_V  => idata_148_pt_V_reg,
      idata_149_pt_V  => idata_149_pt_V_reg,
      idata_150_pt_V  => idata_150_pt_V_reg,
      idata_151_pt_V  => idata_151_pt_V_reg,
      idata_152_pt_V  => idata_152_pt_V_reg,
      idata_153_pt_V  => idata_153_pt_V_reg,
      idata_154_pt_V  => idata_154_pt_V_reg,
      idata_155_pt_V  => idata_155_pt_V_reg,
      idata_156_pt_V  => idata_156_pt_V_reg,
      idata_157_pt_V  => idata_157_pt_V_reg,
      idata_158_pt_V  => idata_158_pt_V_reg,
      idata_159_pt_V  => idata_159_pt_V_reg,
      idata_160_pt_V  => idata_160_pt_V_reg,
      idata_161_pt_V  => idata_161_pt_V_reg,
      idata_162_pt_V  => idata_162_pt_V_reg,
      idata_163_pt_V  => idata_163_pt_V_reg,
      idata_164_pt_V  => idata_164_pt_V_reg,
      idata_165_pt_V  => idata_165_pt_V_reg,
      idata_166_pt_V  => idata_166_pt_V_reg,
      idata_167_pt_V  => idata_167_pt_V_reg,
      idata_168_pt_V  => idata_168_pt_V_reg,
      idata_169_pt_V  => idata_169_pt_V_reg,
      idata_170_pt_V  => idata_170_pt_V_reg,
      idata_171_pt_V  => idata_171_pt_V_reg,
      idata_172_pt_V  => idata_172_pt_V_reg,
      idata_173_pt_V  => idata_173_pt_V_reg,
      idata_174_pt_V  => idata_174_pt_V_reg,
      idata_175_pt_V  => idata_175_pt_V_reg,
      idata_176_pt_V  => idata_176_pt_V_reg,
      idata_177_pt_V  => idata_177_pt_V_reg,
      idata_178_pt_V  => idata_178_pt_V_reg,
      idata_179_pt_V  => idata_179_pt_V_reg,
      idata_180_pt_V  => idata_180_pt_V_reg,
      idata_181_pt_V  => idata_181_pt_V_reg,
      idata_182_pt_V  => idata_182_pt_V_reg,
      idata_183_pt_V  => idata_183_pt_V_reg,
      idata_184_pt_V  => idata_184_pt_V_reg,
      idata_185_pt_V  => idata_185_pt_V_reg,
      idata_186_pt_V  => idata_186_pt_V_reg,
      idata_187_pt_V  => idata_187_pt_V_reg,
      idata_188_pt_V  => idata_188_pt_V_reg,
      idata_189_pt_V  => idata_189_pt_V_reg,
      idata_190_pt_V  => idata_190_pt_V_reg,
      idata_191_pt_V  => idata_191_pt_V_reg,
      idata_192_pt_V  => idata_192_pt_V_reg,
      idata_193_pt_V  => idata_193_pt_V_reg,
      idata_194_pt_V  => idata_194_pt_V_reg,
      idata_195_pt_V  => idata_195_pt_V_reg,
      idata_196_pt_V  => idata_196_pt_V_reg,
      idata_197_pt_V  => idata_197_pt_V_reg,
      idata_198_pt_V  => idata_198_pt_V_reg,
      idata_199_pt_V  => idata_199_pt_V_reg,
      idata_200_pt_V  => idata_200_pt_V_reg,
      idata_201_pt_V  => idata_201_pt_V_reg,
      idata_202_pt_V  => idata_202_pt_V_reg,
      idata_203_pt_V  => idata_203_pt_V_reg,
      idata_204_pt_V  => idata_204_pt_V_reg,
      idata_205_pt_V  => idata_205_pt_V_reg,
      idata_206_pt_V  => idata_206_pt_V_reg,
      idata_207_pt_V  => idata_207_pt_V_reg,
      idata_208_pt_V  => idata_208_pt_V_reg,
      idata_209_pt_V  => idata_209_pt_V_reg,
      idata_210_pt_V  => idata_210_pt_V_reg,
      idata_211_pt_V  => idata_211_pt_V_reg,
      idata_212_pt_V  => idata_212_pt_V_reg,
      idata_213_pt_V  => idata_213_pt_V_reg,
      idata_214_pt_V  => idata_214_pt_V_reg,
      idata_215_pt_V  => idata_215_pt_V_reg,
      idata_216_pt_V  => idata_216_pt_V_reg,
      idata_217_pt_V  => idata_217_pt_V_reg,
      idata_218_pt_V  => idata_218_pt_V_reg,
      idata_219_pt_V  => idata_219_pt_V_reg,
      idata_220_pt_V  => idata_220_pt_V_reg,
      idata_221_pt_V  => idata_221_pt_V_reg,
      idata_222_pt_V  => idata_222_pt_V_reg,
      idata_223_pt_V  => idata_223_pt_V_reg,
      idata_224_pt_V  => idata_224_pt_V_reg,
      idata_225_pt_V  => idata_225_pt_V_reg,
      idata_226_pt_V  => idata_226_pt_V_reg,
      idata_227_pt_V  => idata_227_pt_V_reg,
      idata_228_pt_V  => idata_228_pt_V_reg,
      idata_229_pt_V  => idata_229_pt_V_reg,
      idata_230_pt_V  => idata_230_pt_V_reg,
      idata_231_pt_V  => idata_231_pt_V_reg,
      idata_232_pt_V  => idata_232_pt_V_reg,
      idata_233_pt_V  => idata_233_pt_V_reg,
      idata_234_pt_V  => idata_234_pt_V_reg,
      idata_235_pt_V  => idata_235_pt_V_reg,
      idata_236_pt_V  => idata_236_pt_V_reg,
      idata_237_pt_V  => idata_237_pt_V_reg,
      idata_238_pt_V  => idata_238_pt_V_reg,
      idata_239_pt_V  => idata_239_pt_V_reg,
      idata_240_pt_V  => idata_240_pt_V_reg,
      idata_241_pt_V  => idata_241_pt_V_reg,
      idata_242_pt_V  => idata_242_pt_V_reg,
      idata_243_pt_V  => idata_243_pt_V_reg,
      idata_244_pt_V  => idata_244_pt_V_reg,
      idata_245_pt_V  => idata_245_pt_V_reg,
      idata_246_pt_V  => idata_246_pt_V_reg,
      idata_247_pt_V  => idata_247_pt_V_reg,
      idata_248_pt_V  => idata_248_pt_V_reg,
      idata_249_pt_V  => idata_249_pt_V_reg,
      idata_250_pt_V  => idata_250_pt_V_reg,
      idata_251_pt_V  => idata_251_pt_V_reg,
      idata_252_pt_V  => idata_252_pt_V_reg,
      idata_253_pt_V  => idata_253_pt_V_reg,
      idata_254_pt_V  => idata_254_pt_V_reg,
      idata_255_pt_V  => idata_255_pt_V_reg,
      idata_256_pt_V  => idata_256_pt_V_reg,
      idata_257_pt_V  => idata_257_pt_V_reg,
      idata_258_pt_V  => idata_258_pt_V_reg,
      idata_259_pt_V  => idata_259_pt_V_reg,
      idata_260_pt_V  => idata_260_pt_V_reg,
      idata_261_pt_V  => idata_261_pt_V_reg,
      idata_262_pt_V  => idata_262_pt_V_reg,
      idata_263_pt_V  => idata_263_pt_V_reg,
      idata_264_pt_V  => idata_264_pt_V_reg,
      idata_265_pt_V  => idata_265_pt_V_reg,
      idata_266_pt_V  => idata_266_pt_V_reg,
      idata_267_pt_V  => idata_267_pt_V_reg,
      idata_268_pt_V  => idata_268_pt_V_reg,
      idata_269_pt_V  => idata_269_pt_V_reg,
      idata_270_pt_V  => idata_270_pt_V_reg,
      idata_271_pt_V  => idata_271_pt_V_reg,
      idata_272_pt_V  => idata_272_pt_V_reg,
      idata_273_pt_V  => idata_273_pt_V_reg,
      idata_274_pt_V  => idata_274_pt_V_reg,
      idata_275_pt_V  => idata_275_pt_V_reg,
      idata_276_pt_V  => idata_276_pt_V_reg,
      idata_277_pt_V  => idata_277_pt_V_reg,
      idata_278_pt_V  => idata_278_pt_V_reg,
      idata_279_pt_V  => idata_279_pt_V_reg,
      idata_280_pt_V  => idata_280_pt_V_reg,
      idata_281_pt_V  => idata_281_pt_V_reg,
      idata_282_pt_V  => idata_282_pt_V_reg,
      idata_283_pt_V  => idata_283_pt_V_reg,
      idata_284_pt_V  => idata_284_pt_V_reg,
      idata_285_pt_V  => idata_285_pt_V_reg,
      idata_286_pt_V  => idata_286_pt_V_reg,
      idata_287_pt_V  => idata_287_pt_V_reg,
      idata_288_pt_V  => idata_288_pt_V_reg,
      idata_289_pt_V  => idata_289_pt_V_reg,
      idata_290_pt_V  => idata_290_pt_V_reg,
      idata_291_pt_V  => idata_291_pt_V_reg,
      idata_292_pt_V  => idata_292_pt_V_reg,
      idata_293_pt_V  => idata_293_pt_V_reg,
      idata_294_pt_V  => idata_294_pt_V_reg,
      idata_295_pt_V  => idata_295_pt_V_reg,
      idata_296_pt_V  => idata_296_pt_V_reg,
      idata_297_pt_V  => idata_297_pt_V_reg,
      idata_298_pt_V  => idata_298_pt_V_reg,
      idata_299_pt_V  => idata_299_pt_V_reg,
      idata_300_pt_V  => idata_300_pt_V_reg,
      idata_301_pt_V  => idata_301_pt_V_reg,
      idata_302_pt_V  => idata_302_pt_V_reg,
      idata_303_pt_V  => idata_303_pt_V_reg,
      idata_304_pt_V  => idata_304_pt_V_reg,
      idata_305_pt_V  => idata_305_pt_V_reg,
      idata_306_pt_V  => idata_306_pt_V_reg,
      idata_307_pt_V  => idata_307_pt_V_reg,
      idata_308_pt_V  => idata_308_pt_V_reg,
      idata_309_pt_V  => idata_309_pt_V_reg,
      idata_310_pt_V  => idata_310_pt_V_reg,
      idata_311_pt_V  => idata_311_pt_V_reg,
      idata_312_pt_V  => idata_312_pt_V_reg,
      idata_313_pt_V  => idata_313_pt_V_reg,
      idata_314_pt_V  => idata_314_pt_V_reg,
      idata_315_pt_V  => idata_315_pt_V_reg,
      idata_316_pt_V  => idata_316_pt_V_reg,
      idata_317_pt_V  => idata_317_pt_V_reg,
      idata_318_pt_V  => idata_318_pt_V_reg,
      idata_319_pt_V  => idata_319_pt_V_reg,
      idata_320_pt_V  => idata_320_pt_V_reg,
      idata_321_pt_V  => idata_321_pt_V_reg,
      idata_322_pt_V  => idata_322_pt_V_reg,
      idata_323_pt_V  => idata_323_pt_V_reg,
      idata_324_pt_V  => idata_324_pt_V_reg,
      idata_325_pt_V  => idata_325_pt_V_reg,
      idata_326_pt_V  => idata_326_pt_V_reg,
      idata_327_pt_V  => idata_327_pt_V_reg,
      idata_328_pt_V  => idata_328_pt_V_reg,
      idata_329_pt_V  => idata_329_pt_V_reg,
      idata_330_pt_V  => idata_330_pt_V_reg,
      idata_331_pt_V  => idata_331_pt_V_reg,
      idata_332_pt_V  => idata_332_pt_V_reg,
      idata_333_pt_V  => idata_333_pt_V_reg,
      idata_334_pt_V  => idata_334_pt_V_reg,
      idata_335_pt_V  => idata_335_pt_V_reg,
      idata_336_pt_V  => idata_336_pt_V_reg,
      idata_337_pt_V  => idata_337_pt_V_reg,
      idata_338_pt_V  => idata_338_pt_V_reg,
      idata_339_pt_V  => idata_339_pt_V_reg,
      idata_340_pt_V  => idata_340_pt_V_reg,
      idata_341_pt_V  => idata_341_pt_V_reg,
      idata_342_pt_V  => idata_342_pt_V_reg,
      idata_343_pt_V  => idata_343_pt_V_reg,
      idata_344_pt_V  => idata_344_pt_V_reg,
      idata_345_pt_V  => idata_345_pt_V_reg,
      idata_346_pt_V  => idata_346_pt_V_reg,
      idata_347_pt_V  => idata_347_pt_V_reg,
      idata_348_pt_V  => idata_348_pt_V_reg,
      idata_349_pt_V  => idata_349_pt_V_reg,
      idata_350_pt_V  => idata_350_pt_V_reg,
      idata_351_pt_V  => idata_351_pt_V_reg,
      idata_0_roi_V   => idata_0_roi_V_reg,
      idata_1_roi_V   => idata_1_roi_V_reg,
      idata_2_roi_V   => idata_2_roi_V_reg,
      idata_3_roi_V   => idata_3_roi_V_reg,
      idata_4_roi_V   => idata_4_roi_V_reg,
      idata_5_roi_V   => idata_5_roi_V_reg,
      idata_6_roi_V   => idata_6_roi_V_reg,
      idata_7_roi_V   => idata_7_roi_V_reg,
      idata_8_roi_V   => idata_8_roi_V_reg,
      idata_9_roi_V   => idata_9_roi_V_reg,
      idata_10_roi_V  => idata_10_roi_V_reg,
      idata_11_roi_V  => idata_11_roi_V_reg,
      idata_12_roi_V  => idata_12_roi_V_reg,
      idata_13_roi_V  => idata_13_roi_V_reg,
      idata_14_roi_V  => idata_14_roi_V_reg,
      idata_15_roi_V  => idata_15_roi_V_reg,
      idata_16_roi_V  => idata_16_roi_V_reg,
      idata_17_roi_V  => idata_17_roi_V_reg,
      idata_18_roi_V  => idata_18_roi_V_reg,
      idata_19_roi_V  => idata_19_roi_V_reg,
      idata_20_roi_V  => idata_20_roi_V_reg,
      idata_21_roi_V  => idata_21_roi_V_reg,
      idata_22_roi_V  => idata_22_roi_V_reg,
      idata_23_roi_V  => idata_23_roi_V_reg,
      idata_24_roi_V  => idata_24_roi_V_reg,
      idata_25_roi_V  => idata_25_roi_V_reg,
      idata_26_roi_V  => idata_26_roi_V_reg,
      idata_27_roi_V  => idata_27_roi_V_reg,
      idata_28_roi_V  => idata_28_roi_V_reg,
      idata_29_roi_V  => idata_29_roi_V_reg,
      idata_30_roi_V  => idata_30_roi_V_reg,
      idata_31_roi_V  => idata_31_roi_V_reg,
      idata_32_roi_V  => idata_32_roi_V_reg,
      idata_33_roi_V  => idata_33_roi_V_reg,
      idata_34_roi_V  => idata_34_roi_V_reg,
      idata_35_roi_V  => idata_35_roi_V_reg,
      idata_36_roi_V  => idata_36_roi_V_reg,
      idata_37_roi_V  => idata_37_roi_V_reg,
      idata_38_roi_V  => idata_38_roi_V_reg,
      idata_39_roi_V  => idata_39_roi_V_reg,
      idata_40_roi_V  => idata_40_roi_V_reg,
      idata_41_roi_V  => idata_41_roi_V_reg,
      idata_42_roi_V  => idata_42_roi_V_reg,
      idata_43_roi_V  => idata_43_roi_V_reg,
      idata_44_roi_V  => idata_44_roi_V_reg,
      idata_45_roi_V  => idata_45_roi_V_reg,
      idata_46_roi_V  => idata_46_roi_V_reg,
      idata_47_roi_V  => idata_47_roi_V_reg,
      idata_48_roi_V  => idata_48_roi_V_reg,
      idata_49_roi_V  => idata_49_roi_V_reg,
      idata_50_roi_V  => idata_50_roi_V_reg,
      idata_51_roi_V  => idata_51_roi_V_reg,
      idata_52_roi_V  => idata_52_roi_V_reg,
      idata_53_roi_V  => idata_53_roi_V_reg,
      idata_54_roi_V  => idata_54_roi_V_reg,
      idata_55_roi_V  => idata_55_roi_V_reg,
      idata_56_roi_V  => idata_56_roi_V_reg,
      idata_57_roi_V  => idata_57_roi_V_reg,
      idata_58_roi_V  => idata_58_roi_V_reg,
      idata_59_roi_V  => idata_59_roi_V_reg,
      idata_60_roi_V  => idata_60_roi_V_reg,
      idata_61_roi_V  => idata_61_roi_V_reg,
      idata_62_roi_V  => idata_62_roi_V_reg,
      idata_63_roi_V  => idata_63_roi_V_reg,
      idata_64_roi_V  => idata_64_roi_V_reg,
      idata_65_roi_V  => idata_65_roi_V_reg,
      idata_66_roi_V  => idata_66_roi_V_reg,
      idata_67_roi_V  => idata_67_roi_V_reg,
      idata_68_roi_V  => idata_68_roi_V_reg,
      idata_69_roi_V  => idata_69_roi_V_reg,
      idata_70_roi_V  => idata_70_roi_V_reg,
      idata_71_roi_V  => idata_71_roi_V_reg,
      idata_72_roi_V  => idata_72_roi_V_reg,
      idata_73_roi_V  => idata_73_roi_V_reg,
      idata_74_roi_V  => idata_74_roi_V_reg,
      idata_75_roi_V  => idata_75_roi_V_reg,
      idata_76_roi_V  => idata_76_roi_V_reg,
      idata_77_roi_V  => idata_77_roi_V_reg,
      idata_78_roi_V  => idata_78_roi_V_reg,
      idata_79_roi_V  => idata_79_roi_V_reg,
      idata_80_roi_V  => idata_80_roi_V_reg,
      idata_81_roi_V  => idata_81_roi_V_reg,
      idata_82_roi_V  => idata_82_roi_V_reg,
      idata_83_roi_V  => idata_83_roi_V_reg,
      idata_84_roi_V  => idata_84_roi_V_reg,
      idata_85_roi_V  => idata_85_roi_V_reg,
      idata_86_roi_V  => idata_86_roi_V_reg,
      idata_87_roi_V  => idata_87_roi_V_reg,
      idata_88_roi_V  => idata_88_roi_V_reg,
      idata_89_roi_V  => idata_89_roi_V_reg,
      idata_90_roi_V  => idata_90_roi_V_reg,
      idata_91_roi_V  => idata_91_roi_V_reg,
      idata_92_roi_V  => idata_92_roi_V_reg,
      idata_93_roi_V  => idata_93_roi_V_reg,
      idata_94_roi_V  => idata_94_roi_V_reg,
      idata_95_roi_V  => idata_95_roi_V_reg,
      idata_96_roi_V  => idata_96_roi_V_reg,
      idata_97_roi_V  => idata_97_roi_V_reg,
      idata_98_roi_V  => idata_98_roi_V_reg,
      idata_99_roi_V  => idata_99_roi_V_reg,
      idata_100_roi_V => idata_100_roi_V_reg,
      idata_101_roi_V => idata_101_roi_V_reg,
      idata_102_roi_V => idata_102_roi_V_reg,
      idata_103_roi_V => idata_103_roi_V_reg,
      idata_104_roi_V => idata_104_roi_V_reg,
      idata_105_roi_V => idata_105_roi_V_reg,
      idata_106_roi_V => idata_106_roi_V_reg,
      idata_107_roi_V => idata_107_roi_V_reg,
      idata_108_roi_V => idata_108_roi_V_reg,
      idata_109_roi_V => idata_109_roi_V_reg,
      idata_110_roi_V => idata_110_roi_V_reg,
      idata_111_roi_V => idata_111_roi_V_reg,
      idata_112_roi_V => idata_112_roi_V_reg,
      idata_113_roi_V => idata_113_roi_V_reg,
      idata_114_roi_V => idata_114_roi_V_reg,
      idata_115_roi_V => idata_115_roi_V_reg,
      idata_116_roi_V => idata_116_roi_V_reg,
      idata_117_roi_V => idata_117_roi_V_reg,
      idata_118_roi_V => idata_118_roi_V_reg,
      idata_119_roi_V => idata_119_roi_V_reg,
      idata_120_roi_V => idata_120_roi_V_reg,
      idata_121_roi_V => idata_121_roi_V_reg,
      idata_122_roi_V => idata_122_roi_V_reg,
      idata_123_roi_V => idata_123_roi_V_reg,
      idata_124_roi_V => idata_124_roi_V_reg,
      idata_125_roi_V => idata_125_roi_V_reg,
      idata_126_roi_V => idata_126_roi_V_reg,
      idata_127_roi_V => idata_127_roi_V_reg,
      idata_128_roi_V => idata_128_roi_V_reg,
      idata_129_roi_V => idata_129_roi_V_reg,
      idata_130_roi_V => idata_130_roi_V_reg,
      idata_131_roi_V => idata_131_roi_V_reg,
      idata_132_roi_V => idata_132_roi_V_reg,
      idata_133_roi_V => idata_133_roi_V_reg,
      idata_134_roi_V => idata_134_roi_V_reg,
      idata_135_roi_V => idata_135_roi_V_reg,
      idata_136_roi_V => idata_136_roi_V_reg,
      idata_137_roi_V => idata_137_roi_V_reg,
      idata_138_roi_V => idata_138_roi_V_reg,
      idata_139_roi_V => idata_139_roi_V_reg,
      idata_140_roi_V => idata_140_roi_V_reg,
      idata_141_roi_V => idata_141_roi_V_reg,
      idata_142_roi_V => idata_142_roi_V_reg,
      idata_143_roi_V => idata_143_roi_V_reg,
      idata_144_roi_V => idata_144_roi_V_reg,
      idata_145_roi_V => idata_145_roi_V_reg,
      idata_146_roi_V => idata_146_roi_V_reg,
      idata_147_roi_V => idata_147_roi_V_reg,
      idata_148_roi_V => idata_148_roi_V_reg,
      idata_149_roi_V => idata_149_roi_V_reg,
      idata_150_roi_V => idata_150_roi_V_reg,
      idata_151_roi_V => idata_151_roi_V_reg,
      idata_152_roi_V => idata_152_roi_V_reg,
      idata_153_roi_V => idata_153_roi_V_reg,
      idata_154_roi_V => idata_154_roi_V_reg,
      idata_155_roi_V => idata_155_roi_V_reg,
      idata_156_roi_V => idata_156_roi_V_reg,
      idata_157_roi_V => idata_157_roi_V_reg,
      idata_158_roi_V => idata_158_roi_V_reg,
      idata_159_roi_V => idata_159_roi_V_reg,
      idata_160_roi_V => idata_160_roi_V_reg,
      idata_161_roi_V => idata_161_roi_V_reg,
      idata_162_roi_V => idata_162_roi_V_reg,
      idata_163_roi_V => idata_163_roi_V_reg,
      idata_164_roi_V => idata_164_roi_V_reg,
      idata_165_roi_V => idata_165_roi_V_reg,
      idata_166_roi_V => idata_166_roi_V_reg,
      idata_167_roi_V => idata_167_roi_V_reg,
      idata_168_roi_V => idata_168_roi_V_reg,
      idata_169_roi_V => idata_169_roi_V_reg,
      idata_170_roi_V => idata_170_roi_V_reg,
      idata_171_roi_V => idata_171_roi_V_reg,
      idata_172_roi_V => idata_172_roi_V_reg,
      idata_173_roi_V => idata_173_roi_V_reg,
      idata_174_roi_V => idata_174_roi_V_reg,
      idata_175_roi_V => idata_175_roi_V_reg,
      idata_176_roi_V => idata_176_roi_V_reg,
      idata_177_roi_V => idata_177_roi_V_reg,
      idata_178_roi_V => idata_178_roi_V_reg,
      idata_179_roi_V => idata_179_roi_V_reg,
      idata_180_roi_V => idata_180_roi_V_reg,
      idata_181_roi_V => idata_181_roi_V_reg,
      idata_182_roi_V => idata_182_roi_V_reg,
      idata_183_roi_V => idata_183_roi_V_reg,
      idata_184_roi_V => idata_184_roi_V_reg,
      idata_185_roi_V => idata_185_roi_V_reg,
      idata_186_roi_V => idata_186_roi_V_reg,
      idata_187_roi_V => idata_187_roi_V_reg,
      idata_188_roi_V => idata_188_roi_V_reg,
      idata_189_roi_V => idata_189_roi_V_reg,
      idata_190_roi_V => idata_190_roi_V_reg,
      idata_191_roi_V => idata_191_roi_V_reg,
      idata_192_roi_V => idata_192_roi_V_reg,
      idata_193_roi_V => idata_193_roi_V_reg,
      idata_194_roi_V => idata_194_roi_V_reg,
      idata_195_roi_V => idata_195_roi_V_reg,
      idata_196_roi_V => idata_196_roi_V_reg,
      idata_197_roi_V => idata_197_roi_V_reg,
      idata_198_roi_V => idata_198_roi_V_reg,
      idata_199_roi_V => idata_199_roi_V_reg,
      idata_200_roi_V => idata_200_roi_V_reg,
      idata_201_roi_V => idata_201_roi_V_reg,
      idata_202_roi_V => idata_202_roi_V_reg,
      idata_203_roi_V => idata_203_roi_V_reg,
      idata_204_roi_V => idata_204_roi_V_reg,
      idata_205_roi_V => idata_205_roi_V_reg,
      idata_206_roi_V => idata_206_roi_V_reg,
      idata_207_roi_V => idata_207_roi_V_reg,
      idata_208_roi_V => idata_208_roi_V_reg,
      idata_209_roi_V => idata_209_roi_V_reg,
      idata_210_roi_V => idata_210_roi_V_reg,
      idata_211_roi_V => idata_211_roi_V_reg,
      idata_212_roi_V => idata_212_roi_V_reg,
      idata_213_roi_V => idata_213_roi_V_reg,
      idata_214_roi_V => idata_214_roi_V_reg,
      idata_215_roi_V => idata_215_roi_V_reg,
      idata_216_roi_V => idata_216_roi_V_reg,
      idata_217_roi_V => idata_217_roi_V_reg,
      idata_218_roi_V => idata_218_roi_V_reg,
      idata_219_roi_V => idata_219_roi_V_reg,
      idata_220_roi_V => idata_220_roi_V_reg,
      idata_221_roi_V => idata_221_roi_V_reg,
      idata_222_roi_V => idata_222_roi_V_reg,
      idata_223_roi_V => idata_223_roi_V_reg,
      idata_224_roi_V => idata_224_roi_V_reg,
      idata_225_roi_V => idata_225_roi_V_reg,
      idata_226_roi_V => idata_226_roi_V_reg,
      idata_227_roi_V => idata_227_roi_V_reg,
      idata_228_roi_V => idata_228_roi_V_reg,
      idata_229_roi_V => idata_229_roi_V_reg,
      idata_230_roi_V => idata_230_roi_V_reg,
      idata_231_roi_V => idata_231_roi_V_reg,
      idata_232_roi_V => idata_232_roi_V_reg,
      idata_233_roi_V => idata_233_roi_V_reg,
      idata_234_roi_V => idata_234_roi_V_reg,
      idata_235_roi_V => idata_235_roi_V_reg,
      idata_236_roi_V => idata_236_roi_V_reg,
      idata_237_roi_V => idata_237_roi_V_reg,
      idata_238_roi_V => idata_238_roi_V_reg,
      idata_239_roi_V => idata_239_roi_V_reg,
      idata_240_roi_V => idata_240_roi_V_reg,
      idata_241_roi_V => idata_241_roi_V_reg,
      idata_242_roi_V => idata_242_roi_V_reg,
      idata_243_roi_V => idata_243_roi_V_reg,
      idata_244_roi_V => idata_244_roi_V_reg,
      idata_245_roi_V => idata_245_roi_V_reg,
      idata_246_roi_V => idata_246_roi_V_reg,
      idata_247_roi_V => idata_247_roi_V_reg,
      idata_248_roi_V => idata_248_roi_V_reg,
      idata_249_roi_V => idata_249_roi_V_reg,
      idata_250_roi_V => idata_250_roi_V_reg,
      idata_251_roi_V => idata_251_roi_V_reg,
      idata_252_roi_V => idata_252_roi_V_reg,
      idata_253_roi_V => idata_253_roi_V_reg,
      idata_254_roi_V => idata_254_roi_V_reg,
      idata_255_roi_V => idata_255_roi_V_reg,
      idata_256_roi_V => idata_256_roi_V_reg,
      idata_257_roi_V => idata_257_roi_V_reg,
      idata_258_roi_V => idata_258_roi_V_reg,
      idata_259_roi_V => idata_259_roi_V_reg,
      idata_260_roi_V => idata_260_roi_V_reg,
      idata_261_roi_V => idata_261_roi_V_reg,
      idata_262_roi_V => idata_262_roi_V_reg,
      idata_263_roi_V => idata_263_roi_V_reg,
      idata_264_roi_V => idata_264_roi_V_reg,
      idata_265_roi_V => idata_265_roi_V_reg,
      idata_266_roi_V => idata_266_roi_V_reg,
      idata_267_roi_V => idata_267_roi_V_reg,
      idata_268_roi_V => idata_268_roi_V_reg,
      idata_269_roi_V => idata_269_roi_V_reg,
      idata_270_roi_V => idata_270_roi_V_reg,
      idata_271_roi_V => idata_271_roi_V_reg,
      idata_272_roi_V => idata_272_roi_V_reg,
      idata_273_roi_V => idata_273_roi_V_reg,
      idata_274_roi_V => idata_274_roi_V_reg,
      idata_275_roi_V => idata_275_roi_V_reg,
      idata_276_roi_V => idata_276_roi_V_reg,
      idata_277_roi_V => idata_277_roi_V_reg,
      idata_278_roi_V => idata_278_roi_V_reg,
      idata_279_roi_V => idata_279_roi_V_reg,
      idata_280_roi_V => idata_280_roi_V_reg,
      idata_281_roi_V => idata_281_roi_V_reg,
      idata_282_roi_V => idata_282_roi_V_reg,
      idata_283_roi_V => idata_283_roi_V_reg,
      idata_284_roi_V => idata_284_roi_V_reg,
      idata_285_roi_V => idata_285_roi_V_reg,
      idata_286_roi_V => idata_286_roi_V_reg,
      idata_287_roi_V => idata_287_roi_V_reg,
      idata_288_roi_V => idata_288_roi_V_reg,
      idata_289_roi_V => idata_289_roi_V_reg,
      idata_290_roi_V => idata_290_roi_V_reg,
      idata_291_roi_V => idata_291_roi_V_reg,
      idata_292_roi_V => idata_292_roi_V_reg,
      idata_293_roi_V => idata_293_roi_V_reg,
      idata_294_roi_V => idata_294_roi_V_reg,
      idata_295_roi_V => idata_295_roi_V_reg,
      idata_296_roi_V => idata_296_roi_V_reg,
      idata_297_roi_V => idata_297_roi_V_reg,
      idata_298_roi_V => idata_298_roi_V_reg,
      idata_299_roi_V => idata_299_roi_V_reg,
      idata_300_roi_V => idata_300_roi_V_reg,
      idata_301_roi_V => idata_301_roi_V_reg,
      idata_302_roi_V => idata_302_roi_V_reg,
      idata_303_roi_V => idata_303_roi_V_reg,
      idata_304_roi_V => idata_304_roi_V_reg,
      idata_305_roi_V => idata_305_roi_V_reg,
      idata_306_roi_V => idata_306_roi_V_reg,
      idata_307_roi_V => idata_307_roi_V_reg,
      idata_308_roi_V => idata_308_roi_V_reg,
      idata_309_roi_V => idata_309_roi_V_reg,
      idata_310_roi_V => idata_310_roi_V_reg,
      idata_311_roi_V => idata_311_roi_V_reg,
      idata_312_roi_V => idata_312_roi_V_reg,
      idata_313_roi_V => idata_313_roi_V_reg,
      idata_314_roi_V => idata_314_roi_V_reg,
      idata_315_roi_V => idata_315_roi_V_reg,
      idata_316_roi_V => idata_316_roi_V_reg,
      idata_317_roi_V => idata_317_roi_V_reg,
      idata_318_roi_V => idata_318_roi_V_reg,
      idata_319_roi_V => idata_319_roi_V_reg,
      idata_320_roi_V => idata_320_roi_V_reg,
      idata_321_roi_V => idata_321_roi_V_reg,
      idata_322_roi_V => idata_322_roi_V_reg,
      idata_323_roi_V => idata_323_roi_V_reg,
      idata_324_roi_V => idata_324_roi_V_reg,
      idata_325_roi_V => idata_325_roi_V_reg,
      idata_326_roi_V => idata_326_roi_V_reg,
      idata_327_roi_V => idata_327_roi_V_reg,
      idata_328_roi_V => idata_328_roi_V_reg,
      idata_329_roi_V => idata_329_roi_V_reg,
      idata_330_roi_V => idata_330_roi_V_reg,
      idata_331_roi_V => idata_331_roi_V_reg,
      idata_332_roi_V => idata_332_roi_V_reg,
      idata_333_roi_V => idata_333_roi_V_reg,
      idata_334_roi_V => idata_334_roi_V_reg,
      idata_335_roi_V => idata_335_roi_V_reg,
      idata_336_roi_V => idata_336_roi_V_reg,
      idata_337_roi_V => idata_337_roi_V_reg,
      idata_338_roi_V => idata_338_roi_V_reg,
      idata_339_roi_V => idata_339_roi_V_reg,
      idata_340_roi_V => idata_340_roi_V_reg,
      idata_341_roi_V => idata_341_roi_V_reg,
      idata_342_roi_V => idata_342_roi_V_reg,
      idata_343_roi_V => idata_343_roi_V_reg,
      idata_344_roi_V => idata_344_roi_V_reg,
      idata_345_roi_V => idata_345_roi_V_reg,
      idata_346_roi_V => idata_346_roi_V_reg,
      idata_347_roi_V => idata_347_roi_V_reg,
      idata_348_roi_V => idata_348_roi_V_reg,
      idata_349_roi_V => idata_349_roi_V_reg,
      idata_350_roi_V => idata_350_roi_V_reg,
      idata_351_roi_V => idata_351_roi_V_reg,
      idata_0_flg_V   => idata_0_flg_V_reg,
      idata_1_flg_V   => idata_1_flg_V_reg,
      idata_2_flg_V   => idata_2_flg_V_reg,
      idata_3_flg_V   => idata_3_flg_V_reg,
      idata_4_flg_V   => idata_4_flg_V_reg,
      idata_5_flg_V   => idata_5_flg_V_reg,
      idata_6_flg_V   => idata_6_flg_V_reg,
      idata_7_flg_V   => idata_7_flg_V_reg,
      idata_8_flg_V   => idata_8_flg_V_reg,
      idata_9_flg_V   => idata_9_flg_V_reg,
      idata_10_flg_V  => idata_10_flg_V_reg,
      idata_11_flg_V  => idata_11_flg_V_reg,
      idata_12_flg_V  => idata_12_flg_V_reg,
      idata_13_flg_V  => idata_13_flg_V_reg,
      idata_14_flg_V  => idata_14_flg_V_reg,
      idata_15_flg_V  => idata_15_flg_V_reg,
      idata_16_flg_V  => idata_16_flg_V_reg,
      idata_17_flg_V  => idata_17_flg_V_reg,
      idata_18_flg_V  => idata_18_flg_V_reg,
      idata_19_flg_V  => idata_19_flg_V_reg,
      idata_20_flg_V  => idata_20_flg_V_reg,
      idata_21_flg_V  => idata_21_flg_V_reg,
      idata_22_flg_V  => idata_22_flg_V_reg,
      idata_23_flg_V  => idata_23_flg_V_reg,
      idata_24_flg_V  => idata_24_flg_V_reg,
      idata_25_flg_V  => idata_25_flg_V_reg,
      idata_26_flg_V  => idata_26_flg_V_reg,
      idata_27_flg_V  => idata_27_flg_V_reg,
      idata_28_flg_V  => idata_28_flg_V_reg,
      idata_29_flg_V  => idata_29_flg_V_reg,
      idata_30_flg_V  => idata_30_flg_V_reg,
      idata_31_flg_V  => idata_31_flg_V_reg,
      idata_32_flg_V  => idata_32_flg_V_reg,
      idata_33_flg_V  => idata_33_flg_V_reg,
      idata_34_flg_V  => idata_34_flg_V_reg,
      idata_35_flg_V  => idata_35_flg_V_reg,
      idata_36_flg_V  => idata_36_flg_V_reg,
      idata_37_flg_V  => idata_37_flg_V_reg,
      idata_38_flg_V  => idata_38_flg_V_reg,
      idata_39_flg_V  => idata_39_flg_V_reg,
      idata_40_flg_V  => idata_40_flg_V_reg,
      idata_41_flg_V  => idata_41_flg_V_reg,
      idata_42_flg_V  => idata_42_flg_V_reg,
      idata_43_flg_V  => idata_43_flg_V_reg,
      idata_44_flg_V  => idata_44_flg_V_reg,
      idata_45_flg_V  => idata_45_flg_V_reg,
      idata_46_flg_V  => idata_46_flg_V_reg,
      idata_47_flg_V  => idata_47_flg_V_reg,
      idata_48_flg_V  => idata_48_flg_V_reg,
      idata_49_flg_V  => idata_49_flg_V_reg,
      idata_50_flg_V  => idata_50_flg_V_reg,
      idata_51_flg_V  => idata_51_flg_V_reg,
      idata_52_flg_V  => idata_52_flg_V_reg,
      idata_53_flg_V  => idata_53_flg_V_reg,
      idata_54_flg_V  => idata_54_flg_V_reg,
      idata_55_flg_V  => idata_55_flg_V_reg,
      idata_56_flg_V  => idata_56_flg_V_reg,
      idata_57_flg_V  => idata_57_flg_V_reg,
      idata_58_flg_V  => idata_58_flg_V_reg,
      idata_59_flg_V  => idata_59_flg_V_reg,
      idata_60_flg_V  => idata_60_flg_V_reg,
      idata_61_flg_V  => idata_61_flg_V_reg,
      idata_62_flg_V  => idata_62_flg_V_reg,
      idata_63_flg_V  => idata_63_flg_V_reg,
      idata_64_flg_V  => idata_64_flg_V_reg,
      idata_65_flg_V  => idata_65_flg_V_reg,
      idata_66_flg_V  => idata_66_flg_V_reg,
      idata_67_flg_V  => idata_67_flg_V_reg,
      idata_68_flg_V  => idata_68_flg_V_reg,
      idata_69_flg_V  => idata_69_flg_V_reg,
      idata_70_flg_V  => idata_70_flg_V_reg,
      idata_71_flg_V  => idata_71_flg_V_reg,
      idata_72_flg_V  => idata_72_flg_V_reg,
      idata_73_flg_V  => idata_73_flg_V_reg,
      idata_74_flg_V  => idata_74_flg_V_reg,
      idata_75_flg_V  => idata_75_flg_V_reg,
      idata_76_flg_V  => idata_76_flg_V_reg,
      idata_77_flg_V  => idata_77_flg_V_reg,
      idata_78_flg_V  => idata_78_flg_V_reg,
      idata_79_flg_V  => idata_79_flg_V_reg,
      idata_80_flg_V  => idata_80_flg_V_reg,
      idata_81_flg_V  => idata_81_flg_V_reg,
      idata_82_flg_V  => idata_82_flg_V_reg,
      idata_83_flg_V  => idata_83_flg_V_reg,
      idata_84_flg_V  => idata_84_flg_V_reg,
      idata_85_flg_V  => idata_85_flg_V_reg,
      idata_86_flg_V  => idata_86_flg_V_reg,
      idata_87_flg_V  => idata_87_flg_V_reg,
      idata_88_flg_V  => idata_88_flg_V_reg,
      idata_89_flg_V  => idata_89_flg_V_reg,
      idata_90_flg_V  => idata_90_flg_V_reg,
      idata_91_flg_V  => idata_91_flg_V_reg,
      idata_92_flg_V  => idata_92_flg_V_reg,
      idata_93_flg_V  => idata_93_flg_V_reg,
      idata_94_flg_V  => idata_94_flg_V_reg,
      idata_95_flg_V  => idata_95_flg_V_reg,
      idata_96_flg_V  => idata_96_flg_V_reg,
      idata_97_flg_V  => idata_97_flg_V_reg,
      idata_98_flg_V  => idata_98_flg_V_reg,
      idata_99_flg_V  => idata_99_flg_V_reg,
      idata_100_flg_V => idata_100_flg_V_reg,
      idata_101_flg_V => idata_101_flg_V_reg,
      idata_102_flg_V => idata_102_flg_V_reg,
      idata_103_flg_V => idata_103_flg_V_reg,
      idata_104_flg_V => idata_104_flg_V_reg,
      idata_105_flg_V => idata_105_flg_V_reg,
      idata_106_flg_V => idata_106_flg_V_reg,
      idata_107_flg_V => idata_107_flg_V_reg,
      idata_108_flg_V => idata_108_flg_V_reg,
      idata_109_flg_V => idata_109_flg_V_reg,
      idata_110_flg_V => idata_110_flg_V_reg,
      idata_111_flg_V => idata_111_flg_V_reg,
      idata_112_flg_V => idata_112_flg_V_reg,
      idata_113_flg_V => idata_113_flg_V_reg,
      idata_114_flg_V => idata_114_flg_V_reg,
      idata_115_flg_V => idata_115_flg_V_reg,
      idata_116_flg_V => idata_116_flg_V_reg,
      idata_117_flg_V => idata_117_flg_V_reg,
      idata_118_flg_V => idata_118_flg_V_reg,
      idata_119_flg_V => idata_119_flg_V_reg,
      idata_120_flg_V => idata_120_flg_V_reg,
      idata_121_flg_V => idata_121_flg_V_reg,
      idata_122_flg_V => idata_122_flg_V_reg,
      idata_123_flg_V => idata_123_flg_V_reg,
      idata_124_flg_V => idata_124_flg_V_reg,
      idata_125_flg_V => idata_125_flg_V_reg,
      idata_126_flg_V => idata_126_flg_V_reg,
      idata_127_flg_V => idata_127_flg_V_reg,
      idata_128_flg_V => idata_128_flg_V_reg,
      idata_129_flg_V => idata_129_flg_V_reg,
      idata_130_flg_V => idata_130_flg_V_reg,
      idata_131_flg_V => idata_131_flg_V_reg,
      idata_132_flg_V => idata_132_flg_V_reg,
      idata_133_flg_V => idata_133_flg_V_reg,
      idata_134_flg_V => idata_134_flg_V_reg,
      idata_135_flg_V => idata_135_flg_V_reg,
      idata_136_flg_V => idata_136_flg_V_reg,
      idata_137_flg_V => idata_137_flg_V_reg,
      idata_138_flg_V => idata_138_flg_V_reg,
      idata_139_flg_V => idata_139_flg_V_reg,
      idata_140_flg_V => idata_140_flg_V_reg,
      idata_141_flg_V => idata_141_flg_V_reg,
      idata_142_flg_V => idata_142_flg_V_reg,
      idata_143_flg_V => idata_143_flg_V_reg,
      idata_144_flg_V => idata_144_flg_V_reg,
      idata_145_flg_V => idata_145_flg_V_reg,
      idata_146_flg_V => idata_146_flg_V_reg,
      idata_147_flg_V => idata_147_flg_V_reg,
      idata_148_flg_V => idata_148_flg_V_reg,
      idata_149_flg_V => idata_149_flg_V_reg,
      idata_150_flg_V => idata_150_flg_V_reg,
      idata_151_flg_V => idata_151_flg_V_reg,
      idata_152_flg_V => idata_152_flg_V_reg,
      idata_153_flg_V => idata_153_flg_V_reg,
      idata_154_flg_V => idata_154_flg_V_reg,
      idata_155_flg_V => idata_155_flg_V_reg,
      idata_156_flg_V => idata_156_flg_V_reg,
      idata_157_flg_V => idata_157_flg_V_reg,
      idata_158_flg_V => idata_158_flg_V_reg,
      idata_159_flg_V => idata_159_flg_V_reg,
      idata_160_flg_V => idata_160_flg_V_reg,
      idata_161_flg_V => idata_161_flg_V_reg,
      idata_162_flg_V => idata_162_flg_V_reg,
      idata_163_flg_V => idata_163_flg_V_reg,
      idata_164_flg_V => idata_164_flg_V_reg,
      idata_165_flg_V => idata_165_flg_V_reg,
      idata_166_flg_V => idata_166_flg_V_reg,
      idata_167_flg_V => idata_167_flg_V_reg,
      idata_168_flg_V => idata_168_flg_V_reg,
      idata_169_flg_V => idata_169_flg_V_reg,
      idata_170_flg_V => idata_170_flg_V_reg,
      idata_171_flg_V => idata_171_flg_V_reg,
      idata_172_flg_V => idata_172_flg_V_reg,
      idata_173_flg_V => idata_173_flg_V_reg,
      idata_174_flg_V => idata_174_flg_V_reg,
      idata_175_flg_V => idata_175_flg_V_reg,
      idata_176_flg_V => idata_176_flg_V_reg,
      idata_177_flg_V => idata_177_flg_V_reg,
      idata_178_flg_V => idata_178_flg_V_reg,
      idata_179_flg_V => idata_179_flg_V_reg,
      idata_180_flg_V => idata_180_flg_V_reg,
      idata_181_flg_V => idata_181_flg_V_reg,
      idata_182_flg_V => idata_182_flg_V_reg,
      idata_183_flg_V => idata_183_flg_V_reg,
      idata_184_flg_V => idata_184_flg_V_reg,
      idata_185_flg_V => idata_185_flg_V_reg,
      idata_186_flg_V => idata_186_flg_V_reg,
      idata_187_flg_V => idata_187_flg_V_reg,
      idata_188_flg_V => idata_188_flg_V_reg,
      idata_189_flg_V => idata_189_flg_V_reg,
      idata_190_flg_V => idata_190_flg_V_reg,
      idata_191_flg_V => idata_191_flg_V_reg,
      idata_192_flg_V => idata_192_flg_V_reg,
      idata_193_flg_V => idata_193_flg_V_reg,
      idata_194_flg_V => idata_194_flg_V_reg,
      idata_195_flg_V => idata_195_flg_V_reg,
      idata_196_flg_V => idata_196_flg_V_reg,
      idata_197_flg_V => idata_197_flg_V_reg,
      idata_198_flg_V => idata_198_flg_V_reg,
      idata_199_flg_V => idata_199_flg_V_reg,
      idata_200_flg_V => idata_200_flg_V_reg,
      idata_201_flg_V => idata_201_flg_V_reg,
      idata_202_flg_V => idata_202_flg_V_reg,
      idata_203_flg_V => idata_203_flg_V_reg,
      idata_204_flg_V => idata_204_flg_V_reg,
      idata_205_flg_V => idata_205_flg_V_reg,
      idata_206_flg_V => idata_206_flg_V_reg,
      idata_207_flg_V => idata_207_flg_V_reg,
      idata_208_flg_V => idata_208_flg_V_reg,
      idata_209_flg_V => idata_209_flg_V_reg,
      idata_210_flg_V => idata_210_flg_V_reg,
      idata_211_flg_V => idata_211_flg_V_reg,
      idata_212_flg_V => idata_212_flg_V_reg,
      idata_213_flg_V => idata_213_flg_V_reg,
      idata_214_flg_V => idata_214_flg_V_reg,
      idata_215_flg_V => idata_215_flg_V_reg,
      idata_216_flg_V => idata_216_flg_V_reg,
      idata_217_flg_V => idata_217_flg_V_reg,
      idata_218_flg_V => idata_218_flg_V_reg,
      idata_219_flg_V => idata_219_flg_V_reg,
      idata_220_flg_V => idata_220_flg_V_reg,
      idata_221_flg_V => idata_221_flg_V_reg,
      idata_222_flg_V => idata_222_flg_V_reg,
      idata_223_flg_V => idata_223_flg_V_reg,
      idata_224_flg_V => idata_224_flg_V_reg,
      idata_225_flg_V => idata_225_flg_V_reg,
      idata_226_flg_V => idata_226_flg_V_reg,
      idata_227_flg_V => idata_227_flg_V_reg,
      idata_228_flg_V => idata_228_flg_V_reg,
      idata_229_flg_V => idata_229_flg_V_reg,
      idata_230_flg_V => idata_230_flg_V_reg,
      idata_231_flg_V => idata_231_flg_V_reg,
      idata_232_flg_V => idata_232_flg_V_reg,
      idata_233_flg_V => idata_233_flg_V_reg,
      idata_234_flg_V => idata_234_flg_V_reg,
      idata_235_flg_V => idata_235_flg_V_reg,
      idata_236_flg_V => idata_236_flg_V_reg,
      idata_237_flg_V => idata_237_flg_V_reg,
      idata_238_flg_V => idata_238_flg_V_reg,
      idata_239_flg_V => idata_239_flg_V_reg,
      idata_240_flg_V => idata_240_flg_V_reg,
      idata_241_flg_V => idata_241_flg_V_reg,
      idata_242_flg_V => idata_242_flg_V_reg,
      idata_243_flg_V => idata_243_flg_V_reg,
      idata_244_flg_V => idata_244_flg_V_reg,
      idata_245_flg_V => idata_245_flg_V_reg,
      idata_246_flg_V => idata_246_flg_V_reg,
      idata_247_flg_V => idata_247_flg_V_reg,
      idata_248_flg_V => idata_248_flg_V_reg,
      idata_249_flg_V => idata_249_flg_V_reg,
      idata_250_flg_V => idata_250_flg_V_reg,
      idata_251_flg_V => idata_251_flg_V_reg,
      idata_252_flg_V => idata_252_flg_V_reg,
      idata_253_flg_V => idata_253_flg_V_reg,
      idata_254_flg_V => idata_254_flg_V_reg,
      idata_255_flg_V => idata_255_flg_V_reg,
      idata_256_flg_V => idata_256_flg_V_reg,
      idata_257_flg_V => idata_257_flg_V_reg,
      idata_258_flg_V => idata_258_flg_V_reg,
      idata_259_flg_V => idata_259_flg_V_reg,
      idata_260_flg_V => idata_260_flg_V_reg,
      idata_261_flg_V => idata_261_flg_V_reg,
      idata_262_flg_V => idata_262_flg_V_reg,
      idata_263_flg_V => idata_263_flg_V_reg,
      idata_264_flg_V => idata_264_flg_V_reg,
      idata_265_flg_V => idata_265_flg_V_reg,
      idata_266_flg_V => idata_266_flg_V_reg,
      idata_267_flg_V => idata_267_flg_V_reg,
      idata_268_flg_V => idata_268_flg_V_reg,
      idata_269_flg_V => idata_269_flg_V_reg,
      idata_270_flg_V => idata_270_flg_V_reg,
      idata_271_flg_V => idata_271_flg_V_reg,
      idata_272_flg_V => idata_272_flg_V_reg,
      idata_273_flg_V => idata_273_flg_V_reg,
      idata_274_flg_V => idata_274_flg_V_reg,
      idata_275_flg_V => idata_275_flg_V_reg,
      idata_276_flg_V => idata_276_flg_V_reg,
      idata_277_flg_V => idata_277_flg_V_reg,
      idata_278_flg_V => idata_278_flg_V_reg,
      idata_279_flg_V => idata_279_flg_V_reg,
      idata_280_flg_V => idata_280_flg_V_reg,
      idata_281_flg_V => idata_281_flg_V_reg,
      idata_282_flg_V => idata_282_flg_V_reg,
      idata_283_flg_V => idata_283_flg_V_reg,
      idata_284_flg_V => idata_284_flg_V_reg,
      idata_285_flg_V => idata_285_flg_V_reg,
      idata_286_flg_V => idata_286_flg_V_reg,
      idata_287_flg_V => idata_287_flg_V_reg,
      idata_288_flg_V => idata_288_flg_V_reg,
      idata_289_flg_V => idata_289_flg_V_reg,
      idata_290_flg_V => idata_290_flg_V_reg,
      idata_291_flg_V => idata_291_flg_V_reg,
      idata_292_flg_V => idata_292_flg_V_reg,
      idata_293_flg_V => idata_293_flg_V_reg,
      idata_294_flg_V => idata_294_flg_V_reg,
      idata_295_flg_V => idata_295_flg_V_reg,
      idata_296_flg_V => idata_296_flg_V_reg,
      idata_297_flg_V => idata_297_flg_V_reg,
      idata_298_flg_V => idata_298_flg_V_reg,
      idata_299_flg_V => idata_299_flg_V_reg,
      idata_300_flg_V => idata_300_flg_V_reg,
      idata_301_flg_V => idata_301_flg_V_reg,
      idata_302_flg_V => idata_302_flg_V_reg,
      idata_303_flg_V => idata_303_flg_V_reg,
      idata_304_flg_V => idata_304_flg_V_reg,
      idata_305_flg_V => idata_305_flg_V_reg,
      idata_306_flg_V => idata_306_flg_V_reg,
      idata_307_flg_V => idata_307_flg_V_reg,
      idata_308_flg_V => idata_308_flg_V_reg,
      idata_309_flg_V => idata_309_flg_V_reg,
      idata_310_flg_V => idata_310_flg_V_reg,
      idata_311_flg_V => idata_311_flg_V_reg,
      idata_312_flg_V => idata_312_flg_V_reg,
      idata_313_flg_V => idata_313_flg_V_reg,
      idata_314_flg_V => idata_314_flg_V_reg,
      idata_315_flg_V => idata_315_flg_V_reg,
      idata_316_flg_V => idata_316_flg_V_reg,
      idata_317_flg_V => idata_317_flg_V_reg,
      idata_318_flg_V => idata_318_flg_V_reg,
      idata_319_flg_V => idata_319_flg_V_reg,
      idata_320_flg_V => idata_320_flg_V_reg,
      idata_321_flg_V => idata_321_flg_V_reg,
      idata_322_flg_V => idata_322_flg_V_reg,
      idata_323_flg_V => idata_323_flg_V_reg,
      idata_324_flg_V => idata_324_flg_V_reg,
      idata_325_flg_V => idata_325_flg_V_reg,
      idata_326_flg_V => idata_326_flg_V_reg,
      idata_327_flg_V => idata_327_flg_V_reg,
      idata_328_flg_V => idata_328_flg_V_reg,
      idata_329_flg_V => idata_329_flg_V_reg,
      idata_330_flg_V => idata_330_flg_V_reg,
      idata_331_flg_V => idata_331_flg_V_reg,
      idata_332_flg_V => idata_332_flg_V_reg,
      idata_333_flg_V => idata_333_flg_V_reg,
      idata_334_flg_V => idata_334_flg_V_reg,
      idata_335_flg_V => idata_335_flg_V_reg,
      idata_336_flg_V => idata_336_flg_V_reg,
      idata_337_flg_V => idata_337_flg_V_reg,
      idata_338_flg_V => idata_338_flg_V_reg,
      idata_339_flg_V => idata_339_flg_V_reg,
      idata_340_flg_V => idata_340_flg_V_reg,
      idata_341_flg_V => idata_341_flg_V_reg,
      idata_342_flg_V => idata_342_flg_V_reg,
      idata_343_flg_V => idata_343_flg_V_reg,
      idata_344_flg_V => idata_344_flg_V_reg,
      idata_345_flg_V => idata_345_flg_V_reg,
      idata_346_flg_V => idata_346_flg_V_reg,
      idata_347_flg_V => idata_347_flg_V_reg,
      idata_348_flg_V => idata_348_flg_V_reg,
      idata_349_flg_V => idata_349_flg_V_reg,
      idata_350_flg_V => idata_350_flg_V_reg,
      idata_351_flg_V => idata_351_flg_V_reg,
      odata_0_id_V    => odata_0_id_V,
      odata_1_id_V    => odata_1_id_V,
      odata_2_id_V    => odata_2_id_V,
      odata_3_id_V    => odata_3_id_V,
      odata_4_id_V    => odata_4_id_V,
      odata_5_id_V    => odata_5_id_V,
      odata_6_id_V    => odata_6_id_V,
      odata_7_id_V    => odata_7_id_V,
      odata_8_id_V    => odata_8_id_V,
      odata_9_id_V    => odata_9_id_V,
      odata_10_id_V   => odata_10_id_V,
      odata_11_id_V   => odata_11_id_V,
      odata_12_id_V   => odata_12_id_V,
      odata_13_id_V   => odata_13_id_V,
      odata_14_id_V   => odata_14_id_V,
      odata_15_id_V   => odata_15_id_V,
      odata_0_pt_V    => odata_0_pt_V,
      odata_1_pt_V    => odata_1_pt_V,
      odata_2_pt_V    => odata_2_pt_V,
      odata_3_pt_V    => odata_3_pt_V,
      odata_4_pt_V    => odata_4_pt_V,
      odata_5_pt_V    => odata_5_pt_V,
      odata_6_pt_V    => odata_6_pt_V,
      odata_7_pt_V    => odata_7_pt_V,
      odata_8_pt_V    => odata_8_pt_V,
      odata_9_pt_V    => odata_9_pt_V,
      odata_10_pt_V   => odata_10_pt_V,
      odata_11_pt_V   => odata_11_pt_V,
      odata_12_pt_V   => odata_12_pt_V,
      odata_13_pt_V   => odata_13_pt_V,
      odata_14_pt_V   => odata_14_pt_V,
      odata_15_pt_V   => odata_15_pt_V,
      odata_0_roi_V   => odata_0_roi_V,
      odata_1_roi_V   => odata_1_roi_V,
      odata_2_roi_V   => odata_2_roi_V,
      odata_3_roi_V   => odata_3_roi_V,
      odata_4_roi_V   => odata_4_roi_V,
      odata_5_roi_V   => odata_5_roi_V,
      odata_6_roi_V   => odata_6_roi_V,
      odata_7_roi_V   => odata_7_roi_V,
      odata_8_roi_V   => odata_8_roi_V,
      odata_9_roi_V   => odata_9_roi_V,
      odata_10_roi_V  => odata_10_roi_V,
      odata_11_roi_V  => odata_11_roi_V,
      odata_12_roi_V  => odata_12_roi_V,
      odata_13_roi_V  => odata_13_roi_V,
      odata_14_roi_V  => odata_14_roi_V,
      odata_15_roi_V  => odata_15_roi_V,
      odata_0_flg_V   => odata_0_flg_V,
      odata_1_flg_V   => odata_1_flg_V,
      odata_2_flg_V   => odata_2_flg_V,
      odata_3_flg_V   => odata_3_flg_V,
      odata_4_flg_V   => odata_4_flg_V,
      odata_5_flg_V   => odata_5_flg_V,
      odata_6_flg_V   => odata_6_flg_V,
      odata_7_flg_V   => odata_7_flg_V,
      odata_8_flg_V   => odata_8_flg_V,
      odata_9_flg_V   => odata_9_flg_V,
      odata_10_flg_V  => odata_10_flg_V,
      odata_11_flg_V  => odata_11_flg_V,
      odata_12_flg_V  => odata_12_flg_V,
      odata_13_flg_V  => odata_13_flg_V,
      odata_14_flg_V  => odata_14_flg_V,
      odata_15_flg_V  => odata_15_flg_V);




end architecture rtl;
