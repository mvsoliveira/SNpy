library ieee;
use ieee.std_logic_1164.all;
use IEEE.math_real.all;

package csn_pkg is

	constant MUON_NUMBER : integer := 352;
	constant IDX_WIDTH   : integer := integer(ceil(log(real(MUON_NUMBER), real(2))));
	constant PT_WIDTH    : integer := 4;
	constant word_w      : integer := PT_WIDTH + IDX_WIDTH;

	type muon_type is record
		idx : std_logic_vector(IDX_WIDTH - 1 downto 0);
		pt  : std_logic_vector(PT_WIDTH - 1 downto 0);
	end record;

	type muon_a is array (natural range <>) of muon_type;

	type cmp_cfg is record
		a : natural;
		b : natural;
		p : boolean;
		o : boolean;
		r : boolean;
	end record;

	-- has to be array of array instead of (x,y) array because of issues with synplify
	type pair_cmp_cfg is array (natural range <>) of cmp_cfg;
	type cfg_net_t is array (natural range <>) of pair_cmp_cfg;

	--type cfg_net_t is array (natural range <>, natural range <>) of cmp_cfg;
	function get_cfg(I : integer) return cfg_net_t;

	constant empty_cfg : cfg_net_t := (
		((a => 0, b => 1, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False)),
		((a => 0, b => 2, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False)),
		((a => 1, b => 2, p => False, o => False, r => False), (a => 0, b => 3, p => True, o => False, r => False))
	);

end package csn_pkg;

package body csn_pkg is

	function get_cfg(I : integer) return cfg_net_t is
	begin
		case I is
			-- I=4 batcher odd-even mergesort 
			when 4   => return (
					((a => 0, b => 1, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False)),
					((a => 0, b => 2, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 0, b => 3, p => True, o => False, r => False))
				);
			-- I=8 batcher odd-even mergesort
			when 8   => return (
					((a => 0, b => 1, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False), (a => 4, b => 5, p => False, o => False, r => False), (a => 6, b => 7, p => False, o => False, r => False)),
					((a => 0, b => 2, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False), (a => 4, b => 6, p => False, o => False, r => False), (a => 5, b => 7, p => False, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 0, b => 7, p => True, o => False, r => False), (a => 3, b => 4, p => True, o => False, r => False)),
					((a => 0, b => 4, p => False, o => False, r => False), (a => 1, b => 5, p => False, o => False, r => False), (a => 2, b => 6, p => False, o => False, r => False), (a => 3, b => 7, p => False, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 0, b => 7, p => True, o => False, r => False), (a => 1, b => 6, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 0, b => 7, p => True, o => False, r => False))
				);
			-- I=16 David C. Van Voorhis 16-key sorting network
			when 16  => return (
					((a => 0, b => 1, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False), (a => 4, b => 5, p => False, o => False, r => False), (a => 6, b => 7, p => False, o => False, r => False), (a => 8, b => 9, p => False, o => False, r => False), (a => 10, b => 11, p => False, o => False, r => False), (a => 12, b => 13, p => False, o => False, r => False), (a => 14, b => 15, p => False, o => False, r => False)),
					((a => 0, b => 2, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False), (a => 4, b => 6, p => False, o => False, r => False), (a => 5, b => 7, p => False, o => False, r => False), (a => 8, b => 10, p => False, o => False, r => False), (a => 9, b => 11, p => False, o => False, r => False), (a => 12, b => 14, p => False, o => False, r => False), (a => 13, b => 15, p => False, o => False, r => False)),
					((a => 0, b => 4, p => False, o => False, r => False), (a => 1, b => 5, p => False, o => False, r => False), (a => 2, b => 6, p => False, o => False, r => False), (a => 3, b => 7, p => False, o => False, r => False), (a => 8, b => 12, p => False, o => False, r => False), (a => 9, b => 13, p => False, o => False, r => False), (a => 10, b => 14, p => False, o => False, r => False), (a => 11, b => 15, p => False, o => False, r => False)),
					((a => 0, b => 8, p => False, o => False, r => False), (a => 1, b => 9, p => False, o => False, r => False), (a => 2, b => 10, p => False, o => False, r => False), (a => 3, b => 11, p => False, o => False, r => False), (a => 4, b => 12, p => False, o => False, r => False), (a => 5, b => 13, p => False, o => False, r => False), (a => 6, b => 14, p => False, o => False, r => False), (a => 7, b => 15, p => False, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 4, b => 8, p => False, o => False, r => False), (a => 5, b => 10, p => False, o => False, r => False), (a => 6, b => 9, p => False, o => False, r => False), (a => 0, b => 15, p => True, o => False, r => False)),
					((a => 1, b => 4, p => False, o => False, r => False), (a => 2, b => 8, p => False, o => False, r => False), (a => 3, b => 10, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 6, b => 12, p => False, o => False, r => False), (a => 7, b => 13, p => False, o => False, r => False), (a => 11, b => 14, p => False, o => False, r => False), (a => 0, b => 15, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 0, b => 15, p => True, o => False, r => False), (a => 1, b => 14, p => True, o => False, r => False)),
					((a => 3, b => 6, p => False, o => False, r => False), (a => 5, b => 8, p => False, o => False, r => False), (a => 7, b => 10, p => False, o => False, r => False), (a => 9, b => 12, p => False, o => False, r => False), (a => 0, b => 15, p => True, o => False, r => False), (a => 1, b => 14, p => True, o => False, r => False), (a => 2, b => 13, p => True, o => False, r => False), (a => 4, b => 11, p => True, o => False, r => False)),
					((a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 0, b => 15, p => True, o => False, r => False), (a => 1, b => 14, p => True, o => False, r => False), (a => 2, b => 13, p => True, o => False, r => False))
				);
			when 22  => return (
					((a => 0, b => 1, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False), (a => 4, b => 5, p => False, o => False, r => False), (a => 6, b => 7, p => False, o => False, r => False), (a => 8, b => 9, p => False, o => False, r => False), (a => 10, b => 11, p => False, o => False, r => False), (a => 12, b => 13, p => False, o => False, r => False), (a => 14, b => 15, p => False, o => False, r => False), (a => 16, b => 17, p => False, o => False, r => False), (a => 18, b => 19, p => False, o => False, r => False), (a => 20, b => 21, p => False, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False), (a => 0, b => 5, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False)),
					((a => 6, b => 10, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 8, b => 12, p => False, o => False, r => False), (a => 9, b => 13, p => False, o => False, r => False), (a => 14, b => 18, p => False, o => False, r => False), (a => 15, b => 19, p => False, o => False, r => False), (a => 16, b => 20, p => False, o => False, r => False), (a => 17, b => 21, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 1, b => 4, p => False, o => False, r => False), (a => 0, b => 2, p => False, o => False, r => False)),
					((a => 9, b => 17, p => False, o => False, r => False), (a => 7, b => 15, p => False, o => False, r => False), (a => 11, b => 19, p => False, o => False, r => False), (a => 8, b => 16, p => False, o => False, r => False), (a => 3, b => 12, p => False, o => False, r => False), (a => 0, b => 10, p => False, o => False, r => False), (a => 1, b => 18, p => False, o => False, r => False), (a => 5, b => 20, p => False, o => False, r => False), (a => 13, b => 21, p => False, o => False, r => False), (a => 6, b => 14, p => False, o => False, r => False), (a => 2, b => 4, p => False, o => False, r => False)),
					((a => 0, b => 7, p => False, o => False, r => False), (a => 17, b => 20, p => False, o => False, r => False), (a => 3, b => 15, p => False, o => False, r => False), (a => 9, b => 18, p => False, o => False, r => False), (a => 2, b => 11, p => False, o => False, r => False), (a => 4, b => 16, p => False, o => False, r => False), (a => 5, b => 10, p => False, o => False, r => False), (a => 1, b => 8, p => False, o => False, r => False), (a => 12, b => 19, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 6, b => 21, p => True, o => False, r => False)),
					((a => 20, b => 21, p => False, o => False, r => False), (a => 0, b => 6, p => False, o => False, r => False), (a => 3, b => 8, p => False, o => False, r => False), (a => 12, b => 18, p => False, o => False, r => False), (a => 2, b => 13, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 10, b => 15, p => False, o => False, r => False), (a => 4, b => 7, p => False, o => False, r => False), (a => 11, b => 17, p => False, o => False, r => False), (a => 1, b => 19, p => True, o => False, r => False)),
					((a => 16, b => 20, p => False, o => False, r => False), (a => 18, b => 19, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 12, b => 14, p => False, o => False, r => False), (a => 10, b => 11, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 8, b => 13, p => False, o => False, r => False), (a => 4, b => 5, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False), (a => 2, b => 6, p => False, o => False, r => False), (a => 0, b => 21, p => True, o => False, r => False)),
					((a => 19, b => 20, p => False, o => False, r => False), (a => 16, b => 17, p => False, o => False, r => False), (a => 15, b => 18, p => False, o => False, r => False), (a => 11, b => 14, p => False, o => False, r => False), (a => 9, b => 13, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 4, b => 6, p => False, o => False, r => False), (a => 1, b => 2, p => False, o => False, r => False), (a => 0, b => 21, p => True, o => False, r => False)),
					((a => 18, b => 19, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 13, b => 15, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 8, b => 9, p => False, o => False, r => False), (a => 5, b => 10, p => False, o => False, r => False), (a => 6, b => 7, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False), (a => 0, b => 21, p => True, o => False, r => False), (a => 1, b => 20, p => True, o => False, r => False), (a => 4, b => 17, p => True, o => False, r => False)),
					((a => 17, b => 19, p => False, o => False, r => False), (a => 16, b => 18, p => False, o => False, r => False), (a => 14, b => 15, p => False, o => False, r => False), (a => 12, b => 13, p => False, o => False, r => False), (a => 9, b => 11, p => False, o => False, r => False), (a => 8, b => 10, p => False, o => False, r => False), (a => 5, b => 7, p => False, o => False, r => False), (a => 3, b => 6, p => False, o => False, r => False), (a => 2, b => 4, p => False, o => False, r => False), (a => 0, b => 21, p => True, o => False, r => False), (a => 1, b => 20, p => True, o => False, r => False)),
					((a => 17, b => 18, p => False, o => False, r => False), (a => 15, b => 16, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 0, b => 21, p => True, o => False, r => False), (a => 1, b => 20, p => True, o => False, r => False), (a => 2, b => 19, p => True, o => False, r => False)),
					((a => 16, b => 17, p => False, o => False, r => False), (a => 14, b => 15, p => False, o => False, r => False), (a => 12, b => 13, p => False, o => False, r => False), (a => 10, b => 11, p => False, o => False, r => False), (a => 8, b => 9, p => False, o => False, r => False), (a => 6, b => 7, p => False, o => False, r => False), (a => 4, b => 5, p => False, o => False, r => False), (a => 0, b => 21, p => True, o => False, r => False), (a => 1, b => 20, p => True, o => False, r => False), (a => 2, b => 19, p => True, o => False, r => False), (a => 3, b => 18, p => True, o => False, r => False))
				);
			when 352 => return (
					((a => 0, b => 1, p => False, o => False, r => False), (a => 2, b => 3, p => False, o => False, r => False), (a => 4, b => 5, p => False, o => False, r => False), (a => 6, b => 7, p => False, o => False, r => False), (a => 8, b => 9, p => False, o => False, r => False), (a => 10, b => 11, p => False, o => False, r => False), (a => 12, b => 13, p => False, o => False, r => False), (a => 14, b => 15, p => False, o => False, r => False), (a => 16, b => 17, p => False, o => False, r => False), (a => 18, b => 19, p => False, o => False, r => False), (a => 20, b => 21, p => False, o => False, r => False), (a => 22, b => 23, p => False, o => False, r => False), (a => 24, b => 25, p => False, o => False, r => False), (a => 26, b => 27, p => False, o => False, r => False), (a => 28, b => 29, p => False, o => False, r => False), (a => 30, b => 31, p => False, o => False, r => False), (a => 32, b => 33, p => False, o => False, r => False), (a => 34, b => 35, p => False, o => False, r => False), (a => 36, b => 37, p => False, o => False, r => False), (a => 38, b => 39, p => False, o => False, r => False), (a => 40, b => 41, p => False, o => False, r => False), (a => 42, b => 43, p => False, o => False, r => False), (a => 44, b => 45, p => False, o => False, r => False), (a => 46, b => 47, p => False, o => False, r => False), (a => 48, b => 49, p => False, o => False, r => False), (a => 50, b => 51, p => False, o => False, r => False), (a => 52, b => 53, p => False, o => False, r => False), (a => 54, b => 55, p => False, o => False, r => False), (a => 56, b => 57, p => False, o => False, r => False), (a => 58, b => 59, p => False, o => False, r => False), (a => 60, b => 61, p => False, o => False, r => False), (a => 62, b => 63, p => False, o => False, r => False), (a => 64, b => 65, p => False, o => False, r => False), (a => 66, b => 67, p => False, o => False, r => False), (a => 68, b => 69, p => False, o => False, r => False), (a => 70, b => 71, p => False, o => False, r => False), (a => 72, b => 73, p => False, o => False, r => False), (a => 74, b => 75, p => False, o => False, r => False), (a => 76, b => 77, p => False, o => False, r => False), (a => 78, b => 79, p => False, o => False, r => False), (a => 80, b => 81, p => False, o => False, r => False), (a => 82, b => 83, p => False, o => False, r => False), (a => 84, b => 85, p => False, o => False, r => False), (a => 86, b => 87, p => False, o => False, r => False), (a => 88, b => 89, p => False, o => False, r => False), (a => 90, b => 91, p => False, o => False, r => False), (a => 92, b => 93, p => False, o => False, r => False), (a => 94, b => 95, p => False, o => False, r => False), (a => 96, b => 97, p => False, o => False, r => False), (a => 98, b => 99, p => False, o => False, r => False), (a => 100, b => 101, p => False, o => False, r => False), (a => 102, b => 103, p => False, o => False, r => False), (a => 104, b => 105, p => False, o => False, r => False), (a => 106, b => 107, p => False, o => False, r => False), (a => 108, b => 109, p => False, o => False, r => False), (a => 110, b => 111, p => False, o => False, r => False), (a => 112, b => 113, p => False, o => False, r => False), (a => 114, b => 115, p => False, o => False, r => False), (a => 116, b => 117, p => False, o => False, r => False), (a => 118, b => 119, p => False, o => False, r => False), (a => 120, b => 121, p => False, o => False, r => False), (a => 122, b => 123, p => False, o => False, r => False), (a => 124, b => 125, p => False, o => False, r => False), (a => 126, b => 127, p => False, o => False, r => False), (a => 128, b => 129, p => False, o => False, r => False), (a => 130, b => 131, p => False, o => False, r => False), (a => 132, b => 133, p => False, o => False, r => False), (a => 134, b => 135, p => False, o => False, r => False), (a => 136, b => 137, p => False, o => False, r => False), (a => 138, b => 139, p => False, o => False, r => False), (a => 140, b => 141, p => False, o => False, r => False), (a => 142, b => 143, p => False, o => False, r => False), (a => 144, b => 145, p => False, o => False, r => False), (a => 146, b => 147, p => False, o => False, r => False), (a => 148, b => 149, p => False, o => False, r => False), (a => 150, b => 151, p => False, o => False, r => False), (a => 152, b => 153, p => False, o => False, r => False), (a => 154, b => 155, p => False, o => False, r => False), (a => 156, b => 157, p => False, o => False, r => False), (a => 158, b => 159, p => False, o => False, r => False), (a => 160, b => 161, p => False, o => False, r => False), (a => 162, b => 163, p => False, o => False, r => False), (a => 164, b => 165, p => False, o => False, r => False), (a => 166, b => 167, p => False, o => False, r => False), (a => 168, b => 169, p => False, o => False, r => False), (a => 170, b => 171, p => False, o => False, r => False), (a => 172, b => 173, p => False, o => False, r => False), (a => 174, b => 175, p => False, o => False, r => False), (a => 176, b => 177, p => False, o => False, r => False), (a => 178, b => 179, p => False, o => False, r => False), (a => 180, b => 181, p => False, o => False, r => False), (a => 182, b => 183, p => False, o => False, r => False), (a => 184, b => 185, p => False, o => False, r => False), (a => 186, b => 187, p => False, o => False, r => False), (a => 188, b => 189, p => False, o => False, r => False), (a => 190, b => 191, p => False, o => False, r => False), (a => 192, b => 193, p => False, o => False, r => False), (a => 194, b => 195, p => False, o => False, r => False), (a => 196, b => 197, p => False, o => False, r => False), (a => 198, b => 199, p => False, o => False, r => False), (a => 200, b => 201, p => False, o => False, r => False), (a => 202, b => 203, p => False, o => False, r => False), (a => 204, b => 205, p => False, o => False, r => False), (a => 206, b => 207, p => False, o => False, r => False), (a => 208, b => 209, p => False, o => False, r => False), (a => 210, b => 211, p => False, o => False, r => False), (a => 212, b => 213, p => False, o => False, r => False), (a => 214, b => 215, p => False, o => False, r => False), (a => 216, b => 217, p => False, o => False, r => False), (a => 218, b => 219, p => False, o => False, r => False), (a => 220, b => 221, p => False, o => False, r => False), (a => 222, b => 223, p => False, o => False, r => False), (a => 224, b => 225, p => False, o => False, r => False), (a => 226, b => 227, p => False, o => False, r => False), (a => 228, b => 229, p => False, o => False, r => False), (a => 230, b => 231, p => False, o => False, r => False), (a => 232, b => 233, p => False, o => False, r => False), (a => 234, b => 235, p => False, o => False, r => False), (a => 236, b => 237, p => False, o => False, r => False), (a => 238, b => 239, p => False, o => False, r => False), (a => 240, b => 241, p => False, o => False, r => False), (a => 242, b => 243, p => False, o => False, r => False), (a => 244, b => 245, p => False, o => False, r => False), (a => 246, b => 247, p => False, o => False, r => False), (a => 248, b => 249, p => False, o => False, r => False), (a => 250, b => 251, p => False, o => False, r => False), (a => 252, b => 253, p => False, o => False, r => False), (a => 254, b => 255, p => False, o => False, r => False), (a => 256, b => 257, p => False, o => False, r => False), (a => 258, b => 259, p => False, o => False, r => False), (a => 260, b => 261, p => False, o => False, r => False), (a => 262, b => 263, p => False, o => False, r => False), (a => 264, b => 265, p => False, o => False, r => False), (a => 266, b => 267, p => False, o => False, r => False), (a => 268, b => 269, p => False, o => False, r => False), (a => 270, b => 271, p => False, o => False, r => False), (a => 272, b => 273, p => False, o => False, r => False), (a => 274, b => 275, p => False, o => False, r => False), (a => 276, b => 277, p => False, o => False, r => False), (a => 278, b => 279, p => False, o => False, r => False), (a => 280, b => 281, p => False, o => False, r => False), (a => 282, b => 283, p => False, o => False, r => False), (a => 284, b => 285, p => False, o => False, r => False), (a => 286, b => 287, p => False, o => False, r => False), (a => 288, b => 289, p => False, o => False, r => False), (a => 290, b => 291, p => False, o => False, r => False), (a => 292, b => 293, p => False, o => False, r => False), (a => 294, b => 295, p => False, o => False, r => False), (a => 296, b => 297, p => False, o => False, r => False), (a => 298, b => 299, p => False, o => False, r => False), (a => 300, b => 301, p => False, o => False, r => False), (a => 302, b => 303, p => False, o => False, r => False), (a => 304, b => 305, p => False, o => False, r => False), (a => 306, b => 307, p => False, o => False, r => False), (a => 308, b => 309, p => False, o => False, r => False), (a => 310, b => 311, p => False, o => False, r => False), (a => 312, b => 313, p => False, o => False, r => False), (a => 314, b => 315, p => False, o => False, r => False), (a => 316, b => 317, p => False, o => False, r => False), (a => 318, b => 319, p => False, o => False, r => False), (a => 320, b => 321, p => False, o => False, r => False), (a => 322, b => 323, p => False, o => False, r => False), (a => 324, b => 325, p => False, o => False, r => False), (a => 326, b => 327, p => False, o => False, r => False), (a => 328, b => 329, p => False, o => False, r => False), (a => 330, b => 331, p => False, o => False, r => False), (a => 332, b => 333, p => False, o => False, r => False), (a => 334, b => 335, p => False, o => False, r => False), (a => 336, b => 337, p => False, o => False, r => False), (a => 338, b => 339, p => False, o => False, r => False), (a => 340, b => 341, p => False, o => False, r => False), (a => 342, b => 343, p => False, o => False, r => False), (a => 344, b => 345, p => False, o => False, r => False), (a => 346, b => 347, p => False, o => False, r => False), (a => 348, b => 349, p => False, o => False, r => False), (a => 350, b => 351, p => False, o => False, r => False)),
					((a => 0, b => 2, p => False, o => False, r => False), (a => 1, b => 3, p => False, o => False, r => False), (a => 4, b => 6, p => False, o => False, r => False), (a => 5, b => 7, p => False, o => False, r => False), (a => 8, b => 10, p => False, o => False, r => False), (a => 9, b => 11, p => False, o => False, r => False), (a => 12, b => 14, p => False, o => False, r => False), (a => 13, b => 15, p => False, o => False, r => False), (a => 16, b => 18, p => False, o => False, r => False), (a => 17, b => 19, p => False, o => False, r => False), (a => 20, b => 22, p => False, o => False, r => False), (a => 21, b => 23, p => False, o => False, r => False), (a => 24, b => 26, p => False, o => False, r => False), (a => 25, b => 27, p => False, o => False, r => False), (a => 28, b => 30, p => False, o => False, r => False), (a => 29, b => 31, p => False, o => False, r => False), (a => 32, b => 34, p => False, o => False, r => False), (a => 33, b => 35, p => False, o => False, r => False), (a => 36, b => 38, p => False, o => False, r => False), (a => 37, b => 39, p => False, o => False, r => False), (a => 40, b => 42, p => False, o => False, r => False), (a => 41, b => 43, p => False, o => False, r => False), (a => 44, b => 46, p => False, o => False, r => False), (a => 45, b => 47, p => False, o => False, r => False), (a => 48, b => 50, p => False, o => False, r => False), (a => 49, b => 51, p => False, o => False, r => False), (a => 52, b => 54, p => False, o => False, r => False), (a => 53, b => 55, p => False, o => False, r => False), (a => 56, b => 58, p => False, o => False, r => False), (a => 57, b => 59, p => False, o => False, r => False), (a => 60, b => 62, p => False, o => False, r => False), (a => 61, b => 63, p => False, o => False, r => False), (a => 64, b => 66, p => False, o => False, r => False), (a => 65, b => 67, p => False, o => False, r => False), (a => 68, b => 70, p => False, o => False, r => False), (a => 69, b => 71, p => False, o => False, r => False), (a => 72, b => 74, p => False, o => False, r => False), (a => 73, b => 75, p => False, o => False, r => False), (a => 76, b => 78, p => False, o => False, r => False), (a => 77, b => 79, p => False, o => False, r => False), (a => 80, b => 82, p => False, o => False, r => False), (a => 81, b => 83, p => False, o => False, r => False), (a => 84, b => 86, p => False, o => False, r => False), (a => 85, b => 87, p => False, o => False, r => False), (a => 88, b => 90, p => False, o => False, r => False), (a => 89, b => 91, p => False, o => False, r => False), (a => 92, b => 94, p => False, o => False, r => False), (a => 93, b => 95, p => False, o => False, r => False), (a => 96, b => 98, p => False, o => False, r => False), (a => 97, b => 99, p => False, o => False, r => False), (a => 100, b => 102, p => False, o => False, r => False), (a => 101, b => 103, p => False, o => False, r => False), (a => 104, b => 106, p => False, o => False, r => False), (a => 105, b => 107, p => False, o => False, r => False), (a => 108, b => 110, p => False, o => False, r => False), (a => 109, b => 111, p => False, o => False, r => False), (a => 112, b => 114, p => False, o => False, r => False), (a => 113, b => 115, p => False, o => False, r => False), (a => 116, b => 118, p => False, o => False, r => False), (a => 117, b => 119, p => False, o => False, r => False), (a => 120, b => 122, p => False, o => False, r => False), (a => 121, b => 123, p => False, o => False, r => False), (a => 124, b => 126, p => False, o => False, r => False), (a => 125, b => 127, p => False, o => False, r => False), (a => 128, b => 130, p => False, o => False, r => False), (a => 129, b => 131, p => False, o => False, r => False), (a => 132, b => 134, p => False, o => False, r => False), (a => 133, b => 135, p => False, o => False, r => False), (a => 136, b => 138, p => False, o => False, r => False), (a => 137, b => 139, p => False, o => False, r => False), (a => 140, b => 142, p => False, o => False, r => False), (a => 141, b => 143, p => False, o => False, r => False), (a => 144, b => 146, p => False, o => False, r => False), (a => 145, b => 147, p => False, o => False, r => False), (a => 148, b => 150, p => False, o => False, r => False), (a => 149, b => 151, p => False, o => False, r => False), (a => 152, b => 154, p => False, o => False, r => False), (a => 153, b => 155, p => False, o => False, r => False), (a => 156, b => 158, p => False, o => False, r => False), (a => 157, b => 159, p => False, o => False, r => False), (a => 160, b => 162, p => False, o => False, r => False), (a => 161, b => 163, p => False, o => False, r => False), (a => 164, b => 166, p => False, o => False, r => False), (a => 165, b => 167, p => False, o => False, r => False), (a => 168, b => 170, p => False, o => False, r => False), (a => 169, b => 171, p => False, o => False, r => False), (a => 172, b => 174, p => False, o => False, r => False), (a => 173, b => 175, p => False, o => False, r => False), (a => 176, b => 178, p => False, o => False, r => False), (a => 177, b => 179, p => False, o => False, r => False), (a => 180, b => 182, p => False, o => False, r => False), (a => 181, b => 183, p => False, o => False, r => False), (a => 184, b => 186, p => False, o => False, r => False), (a => 185, b => 187, p => False, o => False, r => False), (a => 188, b => 190, p => False, o => False, r => False), (a => 189, b => 191, p => False, o => False, r => False), (a => 192, b => 194, p => False, o => False, r => False), (a => 193, b => 195, p => False, o => False, r => False), (a => 196, b => 198, p => False, o => False, r => False), (a => 197, b => 199, p => False, o => False, r => False), (a => 200, b => 202, p => False, o => False, r => False), (a => 201, b => 203, p => False, o => False, r => False), (a => 204, b => 206, p => False, o => False, r => False), (a => 205, b => 207, p => False, o => False, r => False), (a => 208, b => 210, p => False, o => False, r => False), (a => 209, b => 211, p => False, o => False, r => False), (a => 212, b => 214, p => False, o => False, r => False), (a => 213, b => 215, p => False, o => False, r => False), (a => 216, b => 218, p => False, o => False, r => False), (a => 217, b => 219, p => False, o => False, r => False), (a => 220, b => 222, p => False, o => False, r => False), (a => 221, b => 223, p => False, o => False, r => False), (a => 224, b => 226, p => False, o => False, r => False), (a => 225, b => 227, p => False, o => False, r => False), (a => 228, b => 230, p => False, o => False, r => False), (a => 229, b => 231, p => False, o => False, r => False), (a => 232, b => 234, p => False, o => False, r => False), (a => 233, b => 235, p => False, o => False, r => False), (a => 236, b => 238, p => False, o => False, r => False), (a => 237, b => 239, p => False, o => False, r => False), (a => 240, b => 242, p => False, o => False, r => False), (a => 241, b => 243, p => False, o => False, r => False), (a => 244, b => 246, p => False, o => False, r => False), (a => 245, b => 247, p => False, o => False, r => False), (a => 248, b => 250, p => False, o => False, r => False), (a => 249, b => 251, p => False, o => False, r => False), (a => 252, b => 254, p => False, o => False, r => False), (a => 253, b => 255, p => False, o => False, r => False), (a => 256, b => 258, p => False, o => False, r => False), (a => 257, b => 259, p => False, o => False, r => False), (a => 260, b => 262, p => False, o => False, r => False), (a => 261, b => 263, p => False, o => False, r => False), (a => 264, b => 266, p => False, o => False, r => False), (a => 265, b => 267, p => False, o => False, r => False), (a => 268, b => 270, p => False, o => False, r => False), (a => 269, b => 271, p => False, o => False, r => False), (a => 272, b => 274, p => False, o => False, r => False), (a => 273, b => 275, p => False, o => False, r => False), (a => 276, b => 278, p => False, o => False, r => False), (a => 277, b => 279, p => False, o => False, r => False), (a => 280, b => 282, p => False, o => False, r => False), (a => 281, b => 283, p => False, o => False, r => False), (a => 284, b => 286, p => False, o => False, r => False), (a => 285, b => 287, p => False, o => False, r => False), (a => 288, b => 290, p => False, o => False, r => False), (a => 289, b => 291, p => False, o => False, r => False), (a => 292, b => 294, p => False, o => False, r => False), (a => 293, b => 295, p => False, o => False, r => False), (a => 296, b => 298, p => False, o => False, r => False), (a => 297, b => 299, p => False, o => False, r => False), (a => 300, b => 302, p => False, o => False, r => False), (a => 301, b => 303, p => False, o => False, r => False), (a => 304, b => 306, p => False, o => False, r => False), (a => 305, b => 307, p => False, o => False, r => False), (a => 308, b => 310, p => False, o => False, r => False), (a => 309, b => 311, p => False, o => False, r => False), (a => 312, b => 314, p => False, o => False, r => False), (a => 313, b => 315, p => False, o => False, r => False), (a => 316, b => 318, p => False, o => False, r => False), (a => 317, b => 319, p => False, o => False, r => False), (a => 320, b => 322, p => False, o => False, r => False), (a => 321, b => 323, p => False, o => False, r => False), (a => 324, b => 326, p => False, o => False, r => False), (a => 325, b => 327, p => False, o => False, r => False), (a => 328, b => 330, p => False, o => False, r => False), (a => 329, b => 331, p => False, o => False, r => False), (a => 332, b => 334, p => False, o => False, r => False), (a => 333, b => 335, p => False, o => False, r => False), (a => 336, b => 338, p => False, o => False, r => False), (a => 337, b => 339, p => False, o => False, r => False), (a => 340, b => 342, p => False, o => False, r => False), (a => 341, b => 343, p => False, o => False, r => False), (a => 344, b => 346, p => False, o => False, r => False), (a => 345, b => 347, p => False, o => False, r => False), (a => 348, b => 350, p => False, o => False, r => False), (a => 349, b => 351, p => False, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 0, b => 4, p => False, o => False, r => False), (a => 3, b => 7, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 8, b => 12, p => False, o => False, r => False), (a => 11, b => 15, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 16, b => 20, p => False, o => False, r => False), (a => 19, b => 23, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 24, b => 28, p => False, o => False, r => False), (a => 27, b => 31, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 32, b => 36, p => False, o => False, r => False), (a => 35, b => 39, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 40, b => 44, p => False, o => False, r => False), (a => 43, b => 47, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 48, b => 52, p => False, o => False, r => False), (a => 51, b => 55, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 56, b => 60, p => False, o => False, r => False), (a => 59, b => 63, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 64, b => 68, p => False, o => False, r => False), (a => 67, b => 71, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 72, b => 76, p => False, o => False, r => False), (a => 75, b => 79, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 80, b => 84, p => False, o => False, r => False), (a => 83, b => 87, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 88, b => 92, p => False, o => False, r => False), (a => 91, b => 95, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 96, b => 100, p => False, o => False, r => False), (a => 99, b => 103, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 104, b => 108, p => False, o => False, r => False), (a => 107, b => 111, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 112, b => 116, p => False, o => False, r => False), (a => 115, b => 119, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 120, b => 124, p => False, o => False, r => False), (a => 123, b => 127, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 128, b => 132, p => False, o => False, r => False), (a => 131, b => 135, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 136, b => 140, p => False, o => False, r => False), (a => 139, b => 143, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 144, b => 148, p => False, o => False, r => False), (a => 147, b => 151, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 152, b => 156, p => False, o => False, r => False), (a => 155, b => 159, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 160, b => 164, p => False, o => False, r => False), (a => 163, b => 167, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 168, b => 172, p => False, o => False, r => False), (a => 171, b => 175, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 176, b => 180, p => False, o => False, r => False), (a => 179, b => 183, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 184, b => 188, p => False, o => False, r => False), (a => 187, b => 191, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 192, b => 196, p => False, o => False, r => False), (a => 195, b => 199, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 200, b => 204, p => False, o => False, r => False), (a => 203, b => 207, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 208, b => 212, p => False, o => False, r => False), (a => 211, b => 215, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 216, b => 220, p => False, o => False, r => False), (a => 219, b => 223, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 224, b => 228, p => False, o => False, r => False), (a => 227, b => 231, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 232, b => 236, p => False, o => False, r => False), (a => 235, b => 239, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 240, b => 244, p => False, o => False, r => False), (a => 243, b => 247, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 248, b => 252, p => False, o => False, r => False), (a => 251, b => 255, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 256, b => 260, p => False, o => False, r => False), (a => 259, b => 263, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 264, b => 268, p => False, o => False, r => False), (a => 267, b => 271, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 272, b => 276, p => False, o => False, r => False), (a => 275, b => 279, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 280, b => 284, p => False, o => False, r => False), (a => 283, b => 287, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 288, b => 292, p => False, o => False, r => False), (a => 291, b => 295, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 296, b => 300, p => False, o => False, r => False), (a => 299, b => 303, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 304, b => 308, p => False, o => False, r => False), (a => 307, b => 311, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 312, b => 316, p => False, o => False, r => False), (a => 315, b => 319, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 320, b => 324, p => False, o => False, r => False), (a => 323, b => 327, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 328, b => 332, p => False, o => False, r => False), (a => 331, b => 335, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 336, b => 340, p => False, o => False, r => False), (a => 339, b => 343, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 344, b => 348, p => False, o => False, r => False), (a => 347, b => 351, p => False, o => False, r => False)),
					((a => 2, b => 6, p => False, o => False, r => False), (a => 1, b => 5, p => False, o => False, r => False), (a => 10, b => 14, p => False, o => False, r => False), (a => 9, b => 13, p => False, o => False, r => False), (a => 0, b => 8, p => False, o => False, r => False), (a => 7, b => 15, p => False, o => False, r => False), (a => 18, b => 22, p => False, o => False, r => False), (a => 17, b => 21, p => False, o => False, r => False), (a => 26, b => 30, p => False, o => False, r => False), (a => 25, b => 29, p => False, o => False, r => False), (a => 16, b => 24, p => False, o => False, r => False), (a => 23, b => 31, p => False, o => False, r => False), (a => 34, b => 38, p => False, o => False, r => False), (a => 33, b => 37, p => False, o => False, r => False), (a => 42, b => 46, p => False, o => False, r => False), (a => 41, b => 45, p => False, o => False, r => False), (a => 32, b => 40, p => False, o => False, r => False), (a => 39, b => 47, p => False, o => False, r => False), (a => 50, b => 54, p => False, o => False, r => False), (a => 49, b => 53, p => False, o => False, r => False), (a => 58, b => 62, p => False, o => False, r => False), (a => 57, b => 61, p => False, o => False, r => False), (a => 48, b => 56, p => False, o => False, r => False), (a => 55, b => 63, p => False, o => False, r => False), (a => 66, b => 70, p => False, o => False, r => False), (a => 65, b => 69, p => False, o => False, r => False), (a => 74, b => 78, p => False, o => False, r => False), (a => 73, b => 77, p => False, o => False, r => False), (a => 64, b => 72, p => False, o => False, r => False), (a => 71, b => 79, p => False, o => False, r => False), (a => 82, b => 86, p => False, o => False, r => False), (a => 81, b => 85, p => False, o => False, r => False), (a => 90, b => 94, p => False, o => False, r => False), (a => 89, b => 93, p => False, o => False, r => False), (a => 80, b => 88, p => False, o => False, r => False), (a => 87, b => 95, p => False, o => False, r => False), (a => 98, b => 102, p => False, o => False, r => False), (a => 97, b => 101, p => False, o => False, r => False), (a => 106, b => 110, p => False, o => False, r => False), (a => 105, b => 109, p => False, o => False, r => False), (a => 96, b => 104, p => False, o => False, r => False), (a => 103, b => 111, p => False, o => False, r => False), (a => 114, b => 118, p => False, o => False, r => False), (a => 113, b => 117, p => False, o => False, r => False), (a => 122, b => 126, p => False, o => False, r => False), (a => 121, b => 125, p => False, o => False, r => False), (a => 112, b => 120, p => False, o => False, r => False), (a => 119, b => 127, p => False, o => False, r => False), (a => 130, b => 134, p => False, o => False, r => False), (a => 129, b => 133, p => False, o => False, r => False), (a => 138, b => 142, p => False, o => False, r => False), (a => 137, b => 141, p => False, o => False, r => False), (a => 128, b => 136, p => False, o => False, r => False), (a => 135, b => 143, p => False, o => False, r => False), (a => 146, b => 150, p => False, o => False, r => False), (a => 145, b => 149, p => False, o => False, r => False), (a => 154, b => 158, p => False, o => False, r => False), (a => 153, b => 157, p => False, o => False, r => False), (a => 144, b => 152, p => False, o => False, r => False), (a => 151, b => 159, p => False, o => False, r => False), (a => 162, b => 166, p => False, o => False, r => False), (a => 161, b => 165, p => False, o => False, r => False), (a => 170, b => 174, p => False, o => False, r => False), (a => 169, b => 173, p => False, o => False, r => False), (a => 160, b => 168, p => False, o => False, r => False), (a => 167, b => 175, p => False, o => False, r => False), (a => 178, b => 182, p => False, o => False, r => False), (a => 177, b => 181, p => False, o => False, r => False), (a => 186, b => 190, p => False, o => False, r => False), (a => 185, b => 189, p => False, o => False, r => False), (a => 176, b => 184, p => False, o => False, r => False), (a => 183, b => 191, p => False, o => False, r => False), (a => 194, b => 198, p => False, o => False, r => False), (a => 193, b => 197, p => False, o => False, r => False), (a => 202, b => 206, p => False, o => False, r => False), (a => 201, b => 205, p => False, o => False, r => False), (a => 192, b => 200, p => False, o => False, r => False), (a => 199, b => 207, p => False, o => False, r => False), (a => 210, b => 214, p => False, o => False, r => False), (a => 209, b => 213, p => False, o => False, r => False), (a => 218, b => 222, p => False, o => False, r => False), (a => 217, b => 221, p => False, o => False, r => False), (a => 208, b => 216, p => False, o => False, r => False), (a => 215, b => 223, p => False, o => False, r => False), (a => 226, b => 230, p => False, o => False, r => False), (a => 225, b => 229, p => False, o => False, r => False), (a => 234, b => 238, p => False, o => False, r => False), (a => 233, b => 237, p => False, o => False, r => False), (a => 224, b => 232, p => False, o => False, r => False), (a => 231, b => 239, p => False, o => False, r => False), (a => 242, b => 246, p => False, o => False, r => False), (a => 241, b => 245, p => False, o => False, r => False), (a => 250, b => 254, p => False, o => False, r => False), (a => 249, b => 253, p => False, o => False, r => False), (a => 240, b => 248, p => False, o => False, r => False), (a => 247, b => 255, p => False, o => False, r => False), (a => 258, b => 262, p => False, o => False, r => False), (a => 257, b => 261, p => False, o => False, r => False), (a => 266, b => 270, p => False, o => False, r => False), (a => 265, b => 269, p => False, o => False, r => False), (a => 256, b => 264, p => False, o => False, r => False), (a => 263, b => 271, p => False, o => False, r => False), (a => 274, b => 278, p => False, o => False, r => False), (a => 273, b => 277, p => False, o => False, r => False), (a => 282, b => 286, p => False, o => False, r => False), (a => 281, b => 285, p => False, o => False, r => False), (a => 272, b => 280, p => False, o => False, r => False), (a => 279, b => 287, p => False, o => False, r => False), (a => 290, b => 294, p => False, o => False, r => False), (a => 289, b => 293, p => False, o => False, r => False), (a => 298, b => 302, p => False, o => False, r => False), (a => 297, b => 301, p => False, o => False, r => False), (a => 288, b => 296, p => False, o => False, r => False), (a => 295, b => 303, p => False, o => False, r => False), (a => 306, b => 310, p => False, o => False, r => False), (a => 305, b => 309, p => False, o => False, r => False), (a => 314, b => 318, p => False, o => False, r => False), (a => 313, b => 317, p => False, o => False, r => False), (a => 304, b => 312, p => False, o => False, r => False), (a => 311, b => 319, p => False, o => False, r => False), (a => 322, b => 326, p => False, o => False, r => False), (a => 321, b => 325, p => False, o => False, r => False), (a => 330, b => 334, p => False, o => False, r => False), (a => 329, b => 333, p => False, o => False, r => False), (a => 320, b => 328, p => False, o => False, r => False), (a => 327, b => 335, p => False, o => False, r => False), (a => 338, b => 342, p => False, o => False, r => False), (a => 337, b => 341, p => False, o => False, r => False), (a => 346, b => 350, p => False, o => False, r => False), (a => 345, b => 349, p => False, o => False, r => False), (a => 336, b => 344, p => False, o => False, r => False), (a => 343, b => 351, p => False, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 11, b => 340, p => True, o => False, r => False), (a => 12, b => 339, p => True, o => False, r => False), (a => 19, b => 332, p => True, o => False, r => False), (a => 20, b => 331, p => True, o => False, r => False), (a => 27, b => 324, p => True, o => False, r => False), (a => 28, b => 323, p => True, o => False, r => False), (a => 35, b => 316, p => True, o => False, r => False), (a => 36, b => 315, p => True, o => False, r => False), (a => 43, b => 308, p => True, o => False, r => False), (a => 44, b => 307, p => True, o => False, r => False), (a => 51, b => 300, p => True, o => False, r => False), (a => 52, b => 299, p => True, o => False, r => False), (a => 59, b => 292, p => True, o => False, r => False), (a => 60, b => 291, p => True, o => False, r => False), (a => 67, b => 284, p => True, o => False, r => False), (a => 68, b => 283, p => True, o => False, r => False), (a => 75, b => 276, p => True, o => False, r => False), (a => 76, b => 275, p => True, o => False, r => False), (a => 83, b => 268, p => True, o => False, r => False), (a => 84, b => 267, p => True, o => False, r => False), (a => 91, b => 260, p => True, o => False, r => False), (a => 92, b => 259, p => True, o => False, r => False), (a => 99, b => 252, p => True, o => False, r => False), (a => 100, b => 251, p => True, o => False, r => False), (a => 107, b => 244, p => True, o => False, r => False), (a => 108, b => 243, p => True, o => False, r => False), (a => 115, b => 236, p => True, o => False, r => False), (a => 116, b => 235, p => True, o => False, r => False), (a => 123, b => 228, p => True, o => False, r => False), (a => 124, b => 227, p => True, o => False, r => False), (a => 131, b => 220, p => True, o => False, r => False), (a => 132, b => 219, p => True, o => False, r => False), (a => 139, b => 212, p => True, o => False, r => False), (a => 140, b => 211, p => True, o => False, r => False), (a => 147, b => 204, p => True, o => False, r => False), (a => 148, b => 203, p => True, o => False, r => False), (a => 155, b => 196, p => True, o => False, r => False), (a => 156, b => 195, p => True, o => False, r => False), (a => 163, b => 188, p => True, o => False, r => False), (a => 164, b => 187, p => True, o => False, r => False), (a => 171, b => 180, p => True, o => False, r => False), (a => 172, b => 179, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 0, b => 16, p => False, o => False, r => False), (a => 15, b => 31, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 32, b => 48, p => False, o => False, r => False), (a => 47, b => 63, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 64, b => 80, p => False, o => False, r => False), (a => 79, b => 95, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 96, b => 112, p => False, o => False, r => False), (a => 111, b => 127, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 128, b => 144, p => False, o => False, r => False), (a => 143, b => 159, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 160, b => 176, p => False, o => False, r => False), (a => 175, b => 191, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 192, b => 208, p => False, o => False, r => False), (a => 207, b => 223, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 224, b => 240, p => False, o => False, r => False), (a => 239, b => 255, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 256, b => 272, p => False, o => False, r => False), (a => 271, b => 287, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 288, b => 304, p => False, o => False, r => False), (a => 303, b => 319, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 320, b => 336, p => False, o => False, r => False), (a => 335, b => 351, p => False, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 8, b => 343, p => True, o => False, r => False), (a => 9, b => 342, p => True, o => False, r => False), (a => 14, b => 337, p => True, o => False, r => False), (a => 17, b => 334, p => True, o => False, r => False), (a => 22, b => 329, p => True, o => False, r => False), (a => 23, b => 328, p => True, o => False, r => False), (a => 24, b => 327, p => True, o => False, r => False), (a => 25, b => 326, p => True, o => False, r => False), (a => 30, b => 321, p => True, o => False, r => False), (a => 33, b => 318, p => True, o => False, r => False), (a => 38, b => 313, p => True, o => False, r => False), (a => 39, b => 312, p => True, o => False, r => False), (a => 40, b => 311, p => True, o => False, r => False), (a => 41, b => 310, p => True, o => False, r => False), (a => 46, b => 305, p => True, o => False, r => False), (a => 49, b => 302, p => True, o => False, r => False), (a => 54, b => 297, p => True, o => False, r => False), (a => 55, b => 296, p => True, o => False, r => False), (a => 56, b => 295, p => True, o => False, r => False), (a => 57, b => 294, p => True, o => False, r => False), (a => 62, b => 289, p => True, o => False, r => False), (a => 65, b => 286, p => True, o => False, r => False), (a => 70, b => 281, p => True, o => False, r => False), (a => 71, b => 280, p => True, o => False, r => False), (a => 72, b => 279, p => True, o => False, r => False), (a => 73, b => 278, p => True, o => False, r => False), (a => 78, b => 273, p => True, o => False, r => False), (a => 81, b => 270, p => True, o => False, r => False), (a => 86, b => 265, p => True, o => False, r => False), (a => 87, b => 264, p => True, o => False, r => False), (a => 88, b => 263, p => True, o => False, r => False), (a => 89, b => 262, p => True, o => False, r => False), (a => 94, b => 257, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 102, b => 249, p => True, o => False, r => False), (a => 103, b => 248, p => True, o => False, r => False), (a => 104, b => 247, p => True, o => False, r => False), (a => 105, b => 246, p => True, o => False, r => False), (a => 110, b => 241, p => True, o => False, r => False), (a => 113, b => 238, p => True, o => False, r => False), (a => 118, b => 233, p => True, o => False, r => False), (a => 119, b => 232, p => True, o => False, r => False), (a => 120, b => 231, p => True, o => False, r => False), (a => 121, b => 230, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 129, b => 222, p => True, o => False, r => False), (a => 134, b => 217, p => True, o => False, r => False), (a => 135, b => 216, p => True, o => False, r => False), (a => 136, b => 215, p => True, o => False, r => False), (a => 137, b => 214, p => True, o => False, r => False), (a => 142, b => 209, p => True, o => False, r => False), (a => 145, b => 206, p => True, o => False, r => False), (a => 150, b => 201, p => True, o => False, r => False), (a => 151, b => 200, p => True, o => False, r => False), (a => 152, b => 199, p => True, o => False, r => False), (a => 153, b => 198, p => True, o => False, r => False), (a => 158, b => 193, p => True, o => False, r => False), (a => 161, b => 190, p => True, o => False, r => False), (a => 166, b => 185, p => True, o => False, r => False), (a => 167, b => 184, p => True, o => False, r => False), (a => 168, b => 183, p => True, o => False, r => False), (a => 169, b => 182, p => True, o => False, r => False), (a => 174, b => 177, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 0, b => 32, p => False, o => False, r => False), (a => 31, b => 63, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 64, b => 96, p => False, o => False, r => False), (a => 95, b => 127, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 128, b => 160, p => False, o => False, r => False), (a => 159, b => 191, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 192, b => 224, p => False, o => False, r => False), (a => 223, b => 255, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 256, b => 288, p => False, o => False, r => False), (a => 287, b => 319, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 7, b => 351, p => True, o => False, r => False), (a => 8, b => 344, p => True, o => False, r => False), (a => 15, b => 343, p => True, o => False, r => False), (a => 16, b => 336, p => True, o => False, r => False), (a => 23, b => 335, p => True, o => False, r => False), (a => 24, b => 328, p => True, o => False, r => False), (a => 39, b => 327, p => True, o => False, r => False), (a => 40, b => 320, p => True, o => False, r => False), (a => 47, b => 312, p => True, o => False, r => False), (a => 48, b => 311, p => True, o => False, r => False), (a => 55, b => 304, p => True, o => False, r => False), (a => 56, b => 303, p => True, o => False, r => False), (a => 71, b => 296, p => True, o => False, r => False), (a => 72, b => 295, p => True, o => False, r => False), (a => 79, b => 280, p => True, o => False, r => False), (a => 80, b => 279, p => True, o => False, r => False), (a => 87, b => 272, p => True, o => False, r => False), (a => 88, b => 271, p => True, o => False, r => False), (a => 103, b => 264, p => True, o => False, r => False), (a => 104, b => 263, p => True, o => False, r => False), (a => 111, b => 248, p => True, o => False, r => False), (a => 112, b => 247, p => True, o => False, r => False), (a => 119, b => 240, p => True, o => False, r => False), (a => 120, b => 239, p => True, o => False, r => False), (a => 135, b => 232, p => True, o => False, r => False), (a => 136, b => 231, p => True, o => False, r => False), (a => 143, b => 216, p => True, o => False, r => False), (a => 144, b => 215, p => True, o => False, r => False), (a => 151, b => 208, p => True, o => False, r => False), (a => 152, b => 207, p => True, o => False, r => False), (a => 167, b => 200, p => True, o => False, r => False), (a => 168, b => 199, p => True, o => False, r => False), (a => 175, b => 184, p => True, o => False, r => False), (a => 176, b => 183, p => True, o => False, r => False)),
					((a => 4, b => 12, p => False, o => False, r => False), (a => 2, b => 10, p => False, o => False, r => False), (a => 6, b => 14, p => False, o => False, r => False), (a => 1, b => 9, p => False, o => False, r => False), (a => 5, b => 13, p => False, o => False, r => False), (a => 3, b => 11, p => False, o => False, r => False), (a => 20, b => 28, p => False, o => False, r => False), (a => 18, b => 26, p => False, o => False, r => False), (a => 22, b => 30, p => False, o => False, r => False), (a => 17, b => 25, p => False, o => False, r => False), (a => 21, b => 29, p => False, o => False, r => False), (a => 19, b => 27, p => False, o => False, r => False), (a => 36, b => 44, p => False, o => False, r => False), (a => 34, b => 42, p => False, o => False, r => False), (a => 38, b => 46, p => False, o => False, r => False), (a => 33, b => 41, p => False, o => False, r => False), (a => 37, b => 45, p => False, o => False, r => False), (a => 35, b => 43, p => False, o => False, r => False), (a => 52, b => 60, p => False, o => False, r => False), (a => 50, b => 58, p => False, o => False, r => False), (a => 54, b => 62, p => False, o => False, r => False), (a => 49, b => 57, p => False, o => False, r => False), (a => 53, b => 61, p => False, o => False, r => False), (a => 51, b => 59, p => False, o => False, r => False), (a => 68, b => 76, p => False, o => False, r => False), (a => 66, b => 74, p => False, o => False, r => False), (a => 70, b => 78, p => False, o => False, r => False), (a => 65, b => 73, p => False, o => False, r => False), (a => 69, b => 77, p => False, o => False, r => False), (a => 67, b => 75, p => False, o => False, r => False), (a => 84, b => 92, p => False, o => False, r => False), (a => 82, b => 90, p => False, o => False, r => False), (a => 86, b => 94, p => False, o => False, r => False), (a => 81, b => 89, p => False, o => False, r => False), (a => 85, b => 93, p => False, o => False, r => False), (a => 83, b => 91, p => False, o => False, r => False), (a => 100, b => 108, p => False, o => False, r => False), (a => 98, b => 106, p => False, o => False, r => False), (a => 102, b => 110, p => False, o => False, r => False), (a => 97, b => 105, p => False, o => False, r => False), (a => 101, b => 109, p => False, o => False, r => False), (a => 99, b => 107, p => False, o => False, r => False), (a => 116, b => 124, p => False, o => False, r => False), (a => 114, b => 122, p => False, o => False, r => False), (a => 118, b => 126, p => False, o => False, r => False), (a => 113, b => 121, p => False, o => False, r => False), (a => 117, b => 125, p => False, o => False, r => False), (a => 115, b => 123, p => False, o => False, r => False), (a => 0, b => 64, p => False, o => False, r => False), (a => 63, b => 127, p => False, o => False, r => False), (a => 132, b => 140, p => False, o => False, r => False), (a => 130, b => 138, p => False, o => False, r => False), (a => 134, b => 142, p => False, o => False, r => False), (a => 129, b => 137, p => False, o => False, r => False), (a => 133, b => 141, p => False, o => False, r => False), (a => 131, b => 139, p => False, o => False, r => False), (a => 148, b => 156, p => False, o => False, r => False), (a => 146, b => 154, p => False, o => False, r => False), (a => 150, b => 158, p => False, o => False, r => False), (a => 145, b => 153, p => False, o => False, r => False), (a => 149, b => 157, p => False, o => False, r => False), (a => 147, b => 155, p => False, o => False, r => False), (a => 164, b => 172, p => False, o => False, r => False), (a => 162, b => 170, p => False, o => False, r => False), (a => 166, b => 174, p => False, o => False, r => False), (a => 161, b => 169, p => False, o => False, r => False), (a => 165, b => 173, p => False, o => False, r => False), (a => 163, b => 171, p => False, o => False, r => False), (a => 180, b => 188, p => False, o => False, r => False), (a => 178, b => 186, p => False, o => False, r => False), (a => 182, b => 190, p => False, o => False, r => False), (a => 177, b => 185, p => False, o => False, r => False), (a => 181, b => 189, p => False, o => False, r => False), (a => 179, b => 187, p => False, o => False, r => False), (a => 196, b => 204, p => False, o => False, r => False), (a => 194, b => 202, p => False, o => False, r => False), (a => 198, b => 206, p => False, o => False, r => False), (a => 193, b => 201, p => False, o => False, r => False), (a => 197, b => 205, p => False, o => False, r => False), (a => 195, b => 203, p => False, o => False, r => False), (a => 212, b => 220, p => False, o => False, r => False), (a => 210, b => 218, p => False, o => False, r => False), (a => 214, b => 222, p => False, o => False, r => False), (a => 209, b => 217, p => False, o => False, r => False), (a => 213, b => 221, p => False, o => False, r => False), (a => 211, b => 219, p => False, o => False, r => False), (a => 228, b => 236, p => False, o => False, r => False), (a => 226, b => 234, p => False, o => False, r => False), (a => 230, b => 238, p => False, o => False, r => False), (a => 225, b => 233, p => False, o => False, r => False), (a => 229, b => 237, p => False, o => False, r => False), (a => 227, b => 235, p => False, o => False, r => False), (a => 244, b => 252, p => False, o => False, r => False), (a => 242, b => 250, p => False, o => False, r => False), (a => 246, b => 254, p => False, o => False, r => False), (a => 241, b => 249, p => False, o => False, r => False), (a => 245, b => 253, p => False, o => False, r => False), (a => 243, b => 251, p => False, o => False, r => False), (a => 128, b => 192, p => False, o => False, r => False), (a => 191, b => 255, p => False, o => False, r => False), (a => 260, b => 268, p => False, o => False, r => False), (a => 258, b => 266, p => False, o => False, r => False), (a => 262, b => 270, p => False, o => False, r => False), (a => 257, b => 265, p => False, o => False, r => False), (a => 261, b => 269, p => False, o => False, r => False), (a => 259, b => 267, p => False, o => False, r => False), (a => 276, b => 284, p => False, o => False, r => False), (a => 274, b => 282, p => False, o => False, r => False), (a => 278, b => 286, p => False, o => False, r => False), (a => 273, b => 281, p => False, o => False, r => False), (a => 277, b => 285, p => False, o => False, r => False), (a => 275, b => 283, p => False, o => False, r => False), (a => 292, b => 300, p => False, o => False, r => False), (a => 290, b => 298, p => False, o => False, r => False), (a => 294, b => 302, p => False, o => False, r => False), (a => 289, b => 297, p => False, o => False, r => False), (a => 293, b => 301, p => False, o => False, r => False), (a => 291, b => 299, p => False, o => False, r => False), (a => 308, b => 316, p => False, o => False, r => False), (a => 306, b => 314, p => False, o => False, r => False), (a => 310, b => 318, p => False, o => False, r => False), (a => 305, b => 313, p => False, o => False, r => False), (a => 309, b => 317, p => False, o => False, r => False), (a => 307, b => 315, p => False, o => False, r => False), (a => 324, b => 332, p => False, o => False, r => False), (a => 322, b => 330, p => False, o => False, r => False), (a => 326, b => 334, p => False, o => False, r => False), (a => 321, b => 329, p => False, o => False, r => False), (a => 325, b => 333, p => False, o => False, r => False), (a => 323, b => 331, p => False, o => False, r => False), (a => 340, b => 348, p => False, o => False, r => False), (a => 338, b => 346, p => False, o => False, r => False), (a => 342, b => 350, p => False, o => False, r => False), (a => 337, b => 345, p => False, o => False, r => False), (a => 341, b => 349, p => False, o => False, r => False), (a => 339, b => 347, p => False, o => False, r => False), (a => 256, b => 320, p => False, o => False, r => False), (a => 7, b => 351, p => True, o => False, r => False), (a => 8, b => 344, p => True, o => False, r => False), (a => 15, b => 343, p => True, o => False, r => False), (a => 16, b => 336, p => True, o => False, r => False), (a => 23, b => 335, p => True, o => False, r => False), (a => 24, b => 328, p => True, o => False, r => False), (a => 31, b => 327, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 39, b => 312, p => True, o => False, r => False), (a => 40, b => 311, p => True, o => False, r => False), (a => 47, b => 304, p => True, o => False, r => False), (a => 48, b => 303, p => True, o => False, r => False), (a => 55, b => 296, p => True, o => False, r => False), (a => 56, b => 295, p => True, o => False, r => False), (a => 71, b => 288, p => True, o => False, r => False), (a => 72, b => 287, p => True, o => False, r => False), (a => 79, b => 280, p => True, o => False, r => False), (a => 80, b => 279, p => True, o => False, r => False), (a => 87, b => 272, p => True, o => False, r => False), (a => 88, b => 271, p => True, o => False, r => False), (a => 95, b => 264, p => True, o => False, r => False), (a => 96, b => 263, p => True, o => False, r => False), (a => 103, b => 248, p => True, o => False, r => False), (a => 104, b => 247, p => True, o => False, r => False), (a => 111, b => 240, p => True, o => False, r => False), (a => 112, b => 239, p => True, o => False, r => False), (a => 119, b => 232, p => True, o => False, r => False), (a => 120, b => 231, p => True, o => False, r => False), (a => 135, b => 224, p => True, o => False, r => False), (a => 136, b => 223, p => True, o => False, r => False), (a => 143, b => 216, p => True, o => False, r => False), (a => 144, b => 215, p => True, o => False, r => False), (a => 151, b => 208, p => True, o => False, r => False), (a => 152, b => 207, p => True, o => False, r => False), (a => 159, b => 200, p => True, o => False, r => False), (a => 160, b => 199, p => True, o => False, r => False), (a => 167, b => 184, p => True, o => False, r => False), (a => 168, b => 183, p => True, o => False, r => False), (a => 175, b => 176, p => True, o => False, r => False)),
					((a => 4, b => 8, p => False, o => False, r => False), (a => 6, b => 10, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 20, b => 24, p => False, o => False, r => False), (a => 22, b => 26, p => False, o => False, r => False), (a => 21, b => 25, p => False, o => False, r => False), (a => 23, b => 27, p => False, o => False, r => False), (a => 36, b => 40, p => False, o => False, r => False), (a => 38, b => 42, p => False, o => False, r => False), (a => 37, b => 41, p => False, o => False, r => False), (a => 39, b => 43, p => False, o => False, r => False), (a => 52, b => 56, p => False, o => False, r => False), (a => 54, b => 58, p => False, o => False, r => False), (a => 53, b => 57, p => False, o => False, r => False), (a => 55, b => 59, p => False, o => False, r => False), (a => 68, b => 72, p => False, o => False, r => False), (a => 70, b => 74, p => False, o => False, r => False), (a => 69, b => 73, p => False, o => False, r => False), (a => 71, b => 75, p => False, o => False, r => False), (a => 84, b => 88, p => False, o => False, r => False), (a => 86, b => 90, p => False, o => False, r => False), (a => 85, b => 89, p => False, o => False, r => False), (a => 87, b => 91, p => False, o => False, r => False), (a => 100, b => 104, p => False, o => False, r => False), (a => 102, b => 106, p => False, o => False, r => False), (a => 101, b => 105, p => False, o => False, r => False), (a => 103, b => 107, p => False, o => False, r => False), (a => 116, b => 120, p => False, o => False, r => False), (a => 118, b => 122, p => False, o => False, r => False), (a => 117, b => 121, p => False, o => False, r => False), (a => 119, b => 123, p => False, o => False, r => False), (a => 132, b => 136, p => False, o => False, r => False), (a => 134, b => 138, p => False, o => False, r => False), (a => 133, b => 137, p => False, o => False, r => False), (a => 135, b => 139, p => False, o => False, r => False), (a => 148, b => 152, p => False, o => False, r => False), (a => 150, b => 154, p => False, o => False, r => False), (a => 149, b => 153, p => False, o => False, r => False), (a => 151, b => 155, p => False, o => False, r => False), (a => 164, b => 168, p => False, o => False, r => False), (a => 166, b => 170, p => False, o => False, r => False), (a => 165, b => 169, p => False, o => False, r => False), (a => 167, b => 171, p => False, o => False, r => False), (a => 180, b => 184, p => False, o => False, r => False), (a => 182, b => 186, p => False, o => False, r => False), (a => 181, b => 185, p => False, o => False, r => False), (a => 183, b => 187, p => False, o => False, r => False), (a => 196, b => 200, p => False, o => False, r => False), (a => 198, b => 202, p => False, o => False, r => False), (a => 197, b => 201, p => False, o => False, r => False), (a => 199, b => 203, p => False, o => False, r => False), (a => 212, b => 216, p => False, o => False, r => False), (a => 214, b => 218, p => False, o => False, r => False), (a => 213, b => 217, p => False, o => False, r => False), (a => 215, b => 219, p => False, o => False, r => False), (a => 228, b => 232, p => False, o => False, r => False), (a => 230, b => 234, p => False, o => False, r => False), (a => 229, b => 233, p => False, o => False, r => False), (a => 231, b => 235, p => False, o => False, r => False), (a => 244, b => 248, p => False, o => False, r => False), (a => 246, b => 250, p => False, o => False, r => False), (a => 245, b => 249, p => False, o => False, r => False), (a => 247, b => 251, p => False, o => False, r => False), (a => 0, b => 128, p => False, o => False, r => False), (a => 127, b => 255, p => False, o => False, r => False), (a => 260, b => 264, p => False, o => False, r => False), (a => 262, b => 266, p => False, o => False, r => False), (a => 261, b => 265, p => False, o => False, r => False), (a => 263, b => 267, p => False, o => False, r => False), (a => 276, b => 280, p => False, o => False, r => False), (a => 278, b => 282, p => False, o => False, r => False), (a => 277, b => 281, p => False, o => False, r => False), (a => 279, b => 283, p => False, o => False, r => False), (a => 292, b => 296, p => False, o => False, r => False), (a => 294, b => 298, p => False, o => False, r => False), (a => 293, b => 297, p => False, o => False, r => False), (a => 295, b => 299, p => False, o => False, r => False), (a => 308, b => 312, p => False, o => False, r => False), (a => 310, b => 314, p => False, o => False, r => False), (a => 309, b => 313, p => False, o => False, r => False), (a => 311, b => 315, p => False, o => False, r => False), (a => 324, b => 328, p => False, o => False, r => False), (a => 326, b => 330, p => False, o => False, r => False), (a => 325, b => 329, p => False, o => False, r => False), (a => 327, b => 331, p => False, o => False, r => False), (a => 340, b => 344, p => False, o => False, r => False), (a => 342, b => 346, p => False, o => False, r => False), (a => 341, b => 345, p => False, o => False, r => False), (a => 343, b => 347, p => False, o => False, r => False), (a => 1, b => 351, p => True, o => False, r => False), (a => 2, b => 350, p => True, o => False, r => False), (a => 3, b => 349, p => True, o => False, r => False), (a => 12, b => 348, p => True, o => False, r => False), (a => 13, b => 339, p => True, o => False, r => False), (a => 14, b => 338, p => True, o => False, r => False), (a => 15, b => 337, p => True, o => False, r => False), (a => 16, b => 336, p => True, o => False, r => False), (a => 17, b => 335, p => True, o => False, r => False), (a => 18, b => 334, p => True, o => False, r => False), (a => 19, b => 333, p => True, o => False, r => False), (a => 28, b => 332, p => True, o => False, r => False), (a => 29, b => 323, p => True, o => False, r => False), (a => 30, b => 322, p => True, o => False, r => False), (a => 31, b => 321, p => True, o => False, r => False), (a => 32, b => 320, p => True, o => False, r => False), (a => 33, b => 319, p => True, o => False, r => False), (a => 34, b => 318, p => True, o => False, r => False), (a => 35, b => 317, p => True, o => False, r => False), (a => 44, b => 316, p => True, o => False, r => False), (a => 45, b => 307, p => True, o => False, r => False), (a => 46, b => 306, p => True, o => False, r => False), (a => 47, b => 305, p => True, o => False, r => False), (a => 48, b => 304, p => True, o => False, r => False), (a => 49, b => 303, p => True, o => False, r => False), (a => 50, b => 302, p => True, o => False, r => False), (a => 51, b => 301, p => True, o => False, r => False), (a => 60, b => 300, p => True, o => False, r => False), (a => 61, b => 291, p => True, o => False, r => False), (a => 62, b => 290, p => True, o => False, r => False), (a => 63, b => 289, p => True, o => False, r => False), (a => 64, b => 288, p => True, o => False, r => False), (a => 65, b => 287, p => True, o => False, r => False), (a => 66, b => 286, p => True, o => False, r => False), (a => 67, b => 285, p => True, o => False, r => False), (a => 76, b => 284, p => True, o => False, r => False), (a => 77, b => 275, p => True, o => False, r => False), (a => 78, b => 274, p => True, o => False, r => False), (a => 79, b => 273, p => True, o => False, r => False), (a => 80, b => 272, p => True, o => False, r => False), (a => 81, b => 271, p => True, o => False, r => False), (a => 82, b => 270, p => True, o => False, r => False), (a => 83, b => 269, p => True, o => False, r => False), (a => 92, b => 268, p => True, o => False, r => False), (a => 93, b => 259, p => True, o => False, r => False), (a => 94, b => 258, p => True, o => False, r => False), (a => 95, b => 257, p => True, o => False, r => False), (a => 96, b => 256, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 98, b => 253, p => True, o => False, r => False), (a => 99, b => 252, p => True, o => False, r => False), (a => 108, b => 243, p => True, o => False, r => False), (a => 109, b => 242, p => True, o => False, r => False), (a => 110, b => 241, p => True, o => False, r => False), (a => 111, b => 240, p => True, o => False, r => False), (a => 112, b => 239, p => True, o => False, r => False), (a => 113, b => 238, p => True, o => False, r => False), (a => 114, b => 237, p => True, o => False, r => False), (a => 115, b => 236, p => True, o => False, r => False), (a => 124, b => 227, p => True, o => False, r => False), (a => 125, b => 226, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 129, b => 224, p => True, o => False, r => False), (a => 130, b => 223, p => True, o => False, r => False), (a => 131, b => 222, p => True, o => False, r => False), (a => 140, b => 221, p => True, o => False, r => False), (a => 141, b => 220, p => True, o => False, r => False), (a => 142, b => 211, p => True, o => False, r => False), (a => 143, b => 210, p => True, o => False, r => False), (a => 144, b => 209, p => True, o => False, r => False), (a => 145, b => 208, p => True, o => False, r => False), (a => 146, b => 207, p => True, o => False, r => False), (a => 147, b => 206, p => True, o => False, r => False), (a => 156, b => 205, p => True, o => False, r => False), (a => 157, b => 204, p => True, o => False, r => False), (a => 158, b => 195, p => True, o => False, r => False), (a => 159, b => 194, p => True, o => False, r => False), (a => 160, b => 193, p => True, o => False, r => False), (a => 161, b => 192, p => True, o => False, r => False), (a => 162, b => 191, p => True, o => False, r => False), (a => 163, b => 190, p => True, o => False, r => False), (a => 172, b => 189, p => True, o => False, r => False), (a => 173, b => 188, p => True, o => False, r => False), (a => 174, b => 179, p => True, o => False, r => False), (a => 175, b => 178, p => True, o => False, r => False), (a => 176, b => 177, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 22, b => 24, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 23, b => 25, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 38, b => 40, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 39, b => 41, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 54, b => 56, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 55, b => 57, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 70, b => 72, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 71, b => 73, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 86, b => 88, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 87, b => 89, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 102, b => 104, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 103, b => 105, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 118, b => 120, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 119, b => 121, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 134, b => 136, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 135, b => 137, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 150, b => 152, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 151, b => 153, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 166, b => 168, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 167, b => 169, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 182, b => 184, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 183, b => 185, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 198, b => 200, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 199, b => 201, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 214, b => 216, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 215, b => 217, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 230, b => 232, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 231, b => 233, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 246, b => 248, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 247, b => 249, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 262, b => 264, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 263, b => 265, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 278, b => 280, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 279, b => 281, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 294, b => 296, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 295, b => 297, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 310, b => 312, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 311, b => 313, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 326, b => 328, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 327, b => 329, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 342, b => 344, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 343, b => 345, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 0, b => 256, p => False, o => False, r => False), (a => 1, b => 351, p => True, o => False, r => False), (a => 14, b => 350, p => True, o => False, r => False), (a => 15, b => 337, p => True, o => False, r => False), (a => 16, b => 336, p => True, o => False, r => False), (a => 17, b => 335, p => True, o => False, r => False), (a => 30, b => 334, p => True, o => False, r => False), (a => 31, b => 321, p => True, o => False, r => False), (a => 32, b => 320, p => True, o => False, r => False), (a => 33, b => 319, p => True, o => False, r => False), (a => 46, b => 318, p => True, o => False, r => False), (a => 47, b => 305, p => True, o => False, r => False), (a => 48, b => 304, p => True, o => False, r => False), (a => 49, b => 303, p => True, o => False, r => False), (a => 62, b => 302, p => True, o => False, r => False), (a => 63, b => 289, p => True, o => False, r => False), (a => 64, b => 288, p => True, o => False, r => False), (a => 65, b => 287, p => True, o => False, r => False), (a => 78, b => 286, p => True, o => False, r => False), (a => 79, b => 273, p => True, o => False, r => False), (a => 80, b => 272, p => True, o => False, r => False), (a => 81, b => 271, p => True, o => False, r => False), (a => 94, b => 270, p => True, o => False, r => False), (a => 95, b => 257, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 110, b => 241, p => True, o => False, r => False), (a => 111, b => 240, p => True, o => False, r => False), (a => 112, b => 239, p => True, o => False, r => False), (a => 113, b => 238, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 129, b => 222, p => True, o => False, r => False), (a => 142, b => 209, p => True, o => False, r => False), (a => 143, b => 208, p => True, o => False, r => False), (a => 144, b => 207, p => True, o => False, r => False), (a => 145, b => 206, p => True, o => False, r => False), (a => 158, b => 193, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 161, b => 190, p => True, o => False, r => False), (a => 174, b => 177, p => True, o => False, r => False), (a => 175, b => 176, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 23, b => 24, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 39, b => 40, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 55, b => 56, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 71, b => 72, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 87, b => 88, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 103, b => 104, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 119, b => 120, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 135, b => 136, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 151, b => 152, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 167, b => 168, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 183, b => 184, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 199, b => 200, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 215, b => 216, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 231, b => 232, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 247, b => 248, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 263, b => 264, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 279, b => 280, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 295, b => 296, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 311, b => 312, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 327, b => 328, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 343, b => 344, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 15, b => 336, p => True, o => False, r => False), (a => 16, b => 335, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 47, b => 304, p => True, o => False, r => False), (a => 48, b => 303, p => True, o => False, r => False), (a => 63, b => 288, p => True, o => False, r => False), (a => 64, b => 287, p => True, o => False, r => False), (a => 79, b => 272, p => True, o => False, r => False), (a => 80, b => 271, p => True, o => False, r => False), (a => 95, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 111, b => 240, p => True, o => False, r => False), (a => 112, b => 239, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 143, b => 208, p => True, o => False, r => False), (a => 144, b => 207, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 175, b => 176, p => True, o => False, r => False)),
					((a => 8, b => 24, p => False, o => False, r => False), (a => 4, b => 20, p => False, o => False, r => False), (a => 12, b => 28, p => False, o => False, r => False), (a => 2, b => 18, p => False, o => False, r => False), (a => 10, b => 26, p => False, o => False, r => False), (a => 6, b => 22, p => False, o => False, r => False), (a => 14, b => 30, p => False, o => False, r => False), (a => 1, b => 17, p => False, o => False, r => False), (a => 9, b => 25, p => False, o => False, r => False), (a => 5, b => 21, p => False, o => False, r => False), (a => 13, b => 29, p => False, o => False, r => False), (a => 3, b => 19, p => False, o => False, r => False), (a => 11, b => 27, p => False, o => False, r => False), (a => 7, b => 23, p => False, o => False, r => False), (a => 40, b => 56, p => False, o => False, r => False), (a => 36, b => 52, p => False, o => False, r => False), (a => 44, b => 60, p => False, o => False, r => False), (a => 34, b => 50, p => False, o => False, r => False), (a => 42, b => 58, p => False, o => False, r => False), (a => 38, b => 54, p => False, o => False, r => False), (a => 46, b => 62, p => False, o => False, r => False), (a => 33, b => 49, p => False, o => False, r => False), (a => 41, b => 57, p => False, o => False, r => False), (a => 37, b => 53, p => False, o => False, r => False), (a => 45, b => 61, p => False, o => False, r => False), (a => 35, b => 51, p => False, o => False, r => False), (a => 43, b => 59, p => False, o => False, r => False), (a => 39, b => 55, p => False, o => False, r => False), (a => 72, b => 88, p => False, o => False, r => False), (a => 68, b => 84, p => False, o => False, r => False), (a => 76, b => 92, p => False, o => False, r => False), (a => 66, b => 82, p => False, o => False, r => False), (a => 74, b => 90, p => False, o => False, r => False), (a => 70, b => 86, p => False, o => False, r => False), (a => 78, b => 94, p => False, o => False, r => False), (a => 65, b => 81, p => False, o => False, r => False), (a => 73, b => 89, p => False, o => False, r => False), (a => 69, b => 85, p => False, o => False, r => False), (a => 77, b => 93, p => False, o => False, r => False), (a => 67, b => 83, p => False, o => False, r => False), (a => 75, b => 91, p => False, o => False, r => False), (a => 71, b => 87, p => False, o => False, r => False), (a => 104, b => 120, p => False, o => False, r => False), (a => 100, b => 116, p => False, o => False, r => False), (a => 108, b => 124, p => False, o => False, r => False), (a => 98, b => 114, p => False, o => False, r => False), (a => 106, b => 122, p => False, o => False, r => False), (a => 102, b => 118, p => False, o => False, r => False), (a => 110, b => 126, p => False, o => False, r => False), (a => 97, b => 113, p => False, o => False, r => False), (a => 105, b => 121, p => False, o => False, r => False), (a => 101, b => 117, p => False, o => False, r => False), (a => 109, b => 125, p => False, o => False, r => False), (a => 99, b => 115, p => False, o => False, r => False), (a => 107, b => 123, p => False, o => False, r => False), (a => 103, b => 119, p => False, o => False, r => False), (a => 136, b => 152, p => False, o => False, r => False), (a => 132, b => 148, p => False, o => False, r => False), (a => 140, b => 156, p => False, o => False, r => False), (a => 130, b => 146, p => False, o => False, r => False), (a => 138, b => 154, p => False, o => False, r => False), (a => 134, b => 150, p => False, o => False, r => False), (a => 142, b => 158, p => False, o => False, r => False), (a => 129, b => 145, p => False, o => False, r => False), (a => 137, b => 153, p => False, o => False, r => False), (a => 133, b => 149, p => False, o => False, r => False), (a => 141, b => 157, p => False, o => False, r => False), (a => 131, b => 147, p => False, o => False, r => False), (a => 139, b => 155, p => False, o => False, r => False), (a => 135, b => 151, p => False, o => False, r => False), (a => 168, b => 184, p => False, o => False, r => False), (a => 164, b => 180, p => False, o => False, r => False), (a => 172, b => 188, p => False, o => False, r => False), (a => 162, b => 178, p => False, o => False, r => False), (a => 170, b => 186, p => False, o => False, r => False), (a => 166, b => 182, p => False, o => False, r => False), (a => 174, b => 190, p => False, o => False, r => False), (a => 161, b => 177, p => False, o => False, r => False), (a => 169, b => 185, p => False, o => False, r => False), (a => 165, b => 181, p => False, o => False, r => False), (a => 173, b => 189, p => False, o => False, r => False), (a => 163, b => 179, p => False, o => False, r => False), (a => 171, b => 187, p => False, o => False, r => False), (a => 167, b => 183, p => False, o => False, r => False), (a => 200, b => 216, p => False, o => False, r => False), (a => 196, b => 212, p => False, o => False, r => False), (a => 204, b => 220, p => False, o => False, r => False), (a => 194, b => 210, p => False, o => False, r => False), (a => 202, b => 218, p => False, o => False, r => False), (a => 198, b => 214, p => False, o => False, r => False), (a => 206, b => 222, p => False, o => False, r => False), (a => 193, b => 209, p => False, o => False, r => False), (a => 201, b => 217, p => False, o => False, r => False), (a => 197, b => 213, p => False, o => False, r => False), (a => 205, b => 221, p => False, o => False, r => False), (a => 195, b => 211, p => False, o => False, r => False), (a => 203, b => 219, p => False, o => False, r => False), (a => 199, b => 215, p => False, o => False, r => False), (a => 232, b => 248, p => False, o => False, r => False), (a => 228, b => 244, p => False, o => False, r => False), (a => 236, b => 252, p => False, o => False, r => False), (a => 226, b => 242, p => False, o => False, r => False), (a => 234, b => 250, p => False, o => False, r => False), (a => 230, b => 246, p => False, o => False, r => False), (a => 238, b => 254, p => False, o => False, r => False), (a => 225, b => 241, p => False, o => False, r => False), (a => 233, b => 249, p => False, o => False, r => False), (a => 229, b => 245, p => False, o => False, r => False), (a => 237, b => 253, p => False, o => False, r => False), (a => 227, b => 243, p => False, o => False, r => False), (a => 235, b => 251, p => False, o => False, r => False), (a => 231, b => 247, p => False, o => False, r => False), (a => 264, b => 280, p => False, o => False, r => False), (a => 260, b => 276, p => False, o => False, r => False), (a => 268, b => 284, p => False, o => False, r => False), (a => 258, b => 274, p => False, o => False, r => False), (a => 266, b => 282, p => False, o => False, r => False), (a => 262, b => 278, p => False, o => False, r => False), (a => 270, b => 286, p => False, o => False, r => False), (a => 257, b => 273, p => False, o => False, r => False), (a => 265, b => 281, p => False, o => False, r => False), (a => 261, b => 277, p => False, o => False, r => False), (a => 269, b => 285, p => False, o => False, r => False), (a => 259, b => 275, p => False, o => False, r => False), (a => 267, b => 283, p => False, o => False, r => False), (a => 263, b => 279, p => False, o => False, r => False), (a => 296, b => 312, p => False, o => False, r => False), (a => 292, b => 308, p => False, o => False, r => False), (a => 300, b => 316, p => False, o => False, r => False), (a => 290, b => 306, p => False, o => False, r => False), (a => 298, b => 314, p => False, o => False, r => False), (a => 294, b => 310, p => False, o => False, r => False), (a => 302, b => 318, p => False, o => False, r => False), (a => 289, b => 305, p => False, o => False, r => False), (a => 297, b => 313, p => False, o => False, r => False), (a => 293, b => 309, p => False, o => False, r => False), (a => 301, b => 317, p => False, o => False, r => False), (a => 291, b => 307, p => False, o => False, r => False), (a => 299, b => 315, p => False, o => False, r => False), (a => 295, b => 311, p => False, o => False, r => False), (a => 328, b => 344, p => False, o => False, r => False), (a => 324, b => 340, p => False, o => False, r => False), (a => 332, b => 348, p => False, o => False, r => False), (a => 322, b => 338, p => False, o => False, r => False), (a => 330, b => 346, p => False, o => False, r => False), (a => 326, b => 342, p => False, o => False, r => False), (a => 334, b => 350, p => False, o => False, r => False), (a => 321, b => 337, p => False, o => False, r => False), (a => 329, b => 345, p => False, o => False, r => False), (a => 325, b => 341, p => False, o => False, r => False), (a => 333, b => 349, p => False, o => False, r => False), (a => 323, b => 339, p => False, o => False, r => False), (a => 331, b => 347, p => False, o => False, r => False), (a => 327, b => 343, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 15, b => 336, p => True, o => False, r => False), (a => 16, b => 335, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 47, b => 304, p => True, o => False, r => False), (a => 48, b => 303, p => True, o => False, r => False), (a => 63, b => 288, p => True, o => False, r => False), (a => 64, b => 287, p => True, o => False, r => False), (a => 79, b => 272, p => True, o => False, r => False), (a => 80, b => 271, p => True, o => False, r => False), (a => 95, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 111, b => 240, p => True, o => False, r => False), (a => 112, b => 239, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 143, b => 208, p => True, o => False, r => False), (a => 144, b => 207, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 175, b => 176, p => True, o => False, r => False)),
					((a => 8, b => 16, p => False, o => False, r => False), (a => 12, b => 20, p => False, o => False, r => False), (a => 10, b => 18, p => False, o => False, r => False), (a => 14, b => 22, p => False, o => False, r => False), (a => 9, b => 17, p => False, o => False, r => False), (a => 13, b => 21, p => False, o => False, r => False), (a => 11, b => 19, p => False, o => False, r => False), (a => 15, b => 23, p => False, o => False, r => False), (a => 40, b => 48, p => False, o => False, r => False), (a => 44, b => 52, p => False, o => False, r => False), (a => 42, b => 50, p => False, o => False, r => False), (a => 46, b => 54, p => False, o => False, r => False), (a => 41, b => 49, p => False, o => False, r => False), (a => 45, b => 53, p => False, o => False, r => False), (a => 43, b => 51, p => False, o => False, r => False), (a => 47, b => 55, p => False, o => False, r => False), (a => 72, b => 80, p => False, o => False, r => False), (a => 76, b => 84, p => False, o => False, r => False), (a => 74, b => 82, p => False, o => False, r => False), (a => 78, b => 86, p => False, o => False, r => False), (a => 73, b => 81, p => False, o => False, r => False), (a => 77, b => 85, p => False, o => False, r => False), (a => 75, b => 83, p => False, o => False, r => False), (a => 79, b => 87, p => False, o => False, r => False), (a => 104, b => 112, p => False, o => False, r => False), (a => 108, b => 116, p => False, o => False, r => False), (a => 106, b => 114, p => False, o => False, r => False), (a => 110, b => 118, p => False, o => False, r => False), (a => 105, b => 113, p => False, o => False, r => False), (a => 109, b => 117, p => False, o => False, r => False), (a => 107, b => 115, p => False, o => False, r => False), (a => 111, b => 119, p => False, o => False, r => False), (a => 136, b => 144, p => False, o => False, r => False), (a => 140, b => 148, p => False, o => False, r => False), (a => 138, b => 146, p => False, o => False, r => False), (a => 142, b => 150, p => False, o => False, r => False), (a => 137, b => 145, p => False, o => False, r => False), (a => 141, b => 149, p => False, o => False, r => False), (a => 139, b => 147, p => False, o => False, r => False), (a => 143, b => 151, p => False, o => False, r => False), (a => 168, b => 176, p => False, o => False, r => False), (a => 172, b => 180, p => False, o => False, r => False), (a => 170, b => 178, p => False, o => False, r => False), (a => 174, b => 182, p => False, o => False, r => False), (a => 169, b => 177, p => False, o => False, r => False), (a => 173, b => 181, p => False, o => False, r => False), (a => 171, b => 179, p => False, o => False, r => False), (a => 175, b => 183, p => False, o => False, r => False), (a => 200, b => 208, p => False, o => False, r => False), (a => 204, b => 212, p => False, o => False, r => False), (a => 202, b => 210, p => False, o => False, r => False), (a => 206, b => 214, p => False, o => False, r => False), (a => 201, b => 209, p => False, o => False, r => False), (a => 205, b => 213, p => False, o => False, r => False), (a => 203, b => 211, p => False, o => False, r => False), (a => 207, b => 215, p => False, o => False, r => False), (a => 232, b => 240, p => False, o => False, r => False), (a => 236, b => 244, p => False, o => False, r => False), (a => 234, b => 242, p => False, o => False, r => False), (a => 238, b => 246, p => False, o => False, r => False), (a => 233, b => 241, p => False, o => False, r => False), (a => 237, b => 245, p => False, o => False, r => False), (a => 235, b => 243, p => False, o => False, r => False), (a => 239, b => 247, p => False, o => False, r => False), (a => 264, b => 272, p => False, o => False, r => False), (a => 268, b => 276, p => False, o => False, r => False), (a => 266, b => 274, p => False, o => False, r => False), (a => 270, b => 278, p => False, o => False, r => False), (a => 265, b => 273, p => False, o => False, r => False), (a => 269, b => 277, p => False, o => False, r => False), (a => 267, b => 275, p => False, o => False, r => False), (a => 271, b => 279, p => False, o => False, r => False), (a => 296, b => 304, p => False, o => False, r => False), (a => 300, b => 308, p => False, o => False, r => False), (a => 298, b => 306, p => False, o => False, r => False), (a => 302, b => 310, p => False, o => False, r => False), (a => 297, b => 305, p => False, o => False, r => False), (a => 301, b => 309, p => False, o => False, r => False), (a => 299, b => 307, p => False, o => False, r => False), (a => 303, b => 311, p => False, o => False, r => False), (a => 328, b => 336, p => False, o => False, r => False), (a => 332, b => 340, p => False, o => False, r => False), (a => 330, b => 338, p => False, o => False, r => False), (a => 334, b => 342, p => False, o => False, r => False), (a => 329, b => 337, p => False, o => False, r => False), (a => 333, b => 341, p => False, o => False, r => False), (a => 331, b => 339, p => False, o => False, r => False), (a => 335, b => 343, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 24, b => 327, p => True, o => False, r => False), (a => 25, b => 326, p => True, o => False, r => False), (a => 26, b => 325, p => True, o => False, r => False), (a => 27, b => 324, p => True, o => False, r => False), (a => 28, b => 323, p => True, o => False, r => False), (a => 29, b => 322, p => True, o => False, r => False), (a => 30, b => 321, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 33, b => 318, p => True, o => False, r => False), (a => 34, b => 317, p => True, o => False, r => False), (a => 35, b => 316, p => True, o => False, r => False), (a => 36, b => 315, p => True, o => False, r => False), (a => 37, b => 314, p => True, o => False, r => False), (a => 38, b => 313, p => True, o => False, r => False), (a => 39, b => 312, p => True, o => False, r => False), (a => 56, b => 295, p => True, o => False, r => False), (a => 57, b => 294, p => True, o => False, r => False), (a => 58, b => 293, p => True, o => False, r => False), (a => 59, b => 292, p => True, o => False, r => False), (a => 60, b => 291, p => True, o => False, r => False), (a => 61, b => 290, p => True, o => False, r => False), (a => 62, b => 289, p => True, o => False, r => False), (a => 63, b => 288, p => True, o => False, r => False), (a => 64, b => 287, p => True, o => False, r => False), (a => 65, b => 286, p => True, o => False, r => False), (a => 66, b => 285, p => True, o => False, r => False), (a => 67, b => 284, p => True, o => False, r => False), (a => 68, b => 283, p => True, o => False, r => False), (a => 69, b => 282, p => True, o => False, r => False), (a => 70, b => 281, p => True, o => False, r => False), (a => 71, b => 280, p => True, o => False, r => False), (a => 88, b => 263, p => True, o => False, r => False), (a => 89, b => 262, p => True, o => False, r => False), (a => 90, b => 261, p => True, o => False, r => False), (a => 91, b => 260, p => True, o => False, r => False), (a => 92, b => 259, p => True, o => False, r => False), (a => 93, b => 258, p => True, o => False, r => False), (a => 94, b => 257, p => True, o => False, r => False), (a => 95, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 98, b => 253, p => True, o => False, r => False), (a => 99, b => 252, p => True, o => False, r => False), (a => 100, b => 251, p => True, o => False, r => False), (a => 101, b => 250, p => True, o => False, r => False), (a => 102, b => 249, p => True, o => False, r => False), (a => 103, b => 248, p => True, o => False, r => False), (a => 120, b => 231, p => True, o => False, r => False), (a => 121, b => 230, p => True, o => False, r => False), (a => 122, b => 229, p => True, o => False, r => False), (a => 123, b => 228, p => True, o => False, r => False), (a => 124, b => 227, p => True, o => False, r => False), (a => 125, b => 226, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 129, b => 222, p => True, o => False, r => False), (a => 130, b => 221, p => True, o => False, r => False), (a => 131, b => 220, p => True, o => False, r => False), (a => 132, b => 219, p => True, o => False, r => False), (a => 133, b => 218, p => True, o => False, r => False), (a => 134, b => 217, p => True, o => False, r => False), (a => 135, b => 216, p => True, o => False, r => False), (a => 152, b => 199, p => True, o => False, r => False), (a => 153, b => 198, p => True, o => False, r => False), (a => 154, b => 197, p => True, o => False, r => False), (a => 155, b => 196, p => True, o => False, r => False), (a => 156, b => 195, p => True, o => False, r => False), (a => 157, b => 194, p => True, o => False, r => False), (a => 158, b => 193, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 161, b => 190, p => True, o => False, r => False), (a => 162, b => 189, p => True, o => False, r => False), (a => 163, b => 188, p => True, o => False, r => False), (a => 164, b => 187, p => True, o => False, r => False), (a => 165, b => 186, p => True, o => False, r => False), (a => 166, b => 185, p => True, o => False, r => False), (a => 167, b => 184, p => True, o => False, r => False)),
					((a => 4, b => 8, p => False, o => False, r => False), (a => 12, b => 16, p => False, o => False, r => False), (a => 20, b => 24, p => False, o => False, r => False), (a => 6, b => 10, p => False, o => False, r => False), (a => 14, b => 18, p => False, o => False, r => False), (a => 22, b => 26, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 13, b => 17, p => False, o => False, r => False), (a => 21, b => 25, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 15, b => 19, p => False, o => False, r => False), (a => 23, b => 27, p => False, o => False, r => False), (a => 36, b => 40, p => False, o => False, r => False), (a => 44, b => 48, p => False, o => False, r => False), (a => 52, b => 56, p => False, o => False, r => False), (a => 38, b => 42, p => False, o => False, r => False), (a => 46, b => 50, p => False, o => False, r => False), (a => 54, b => 58, p => False, o => False, r => False), (a => 37, b => 41, p => False, o => False, r => False), (a => 45, b => 49, p => False, o => False, r => False), (a => 53, b => 57, p => False, o => False, r => False), (a => 39, b => 43, p => False, o => False, r => False), (a => 47, b => 51, p => False, o => False, r => False), (a => 55, b => 59, p => False, o => False, r => False), (a => 68, b => 72, p => False, o => False, r => False), (a => 76, b => 80, p => False, o => False, r => False), (a => 84, b => 88, p => False, o => False, r => False), (a => 70, b => 74, p => False, o => False, r => False), (a => 78, b => 82, p => False, o => False, r => False), (a => 86, b => 90, p => False, o => False, r => False), (a => 69, b => 73, p => False, o => False, r => False), (a => 77, b => 81, p => False, o => False, r => False), (a => 85, b => 89, p => False, o => False, r => False), (a => 71, b => 75, p => False, o => False, r => False), (a => 79, b => 83, p => False, o => False, r => False), (a => 87, b => 91, p => False, o => False, r => False), (a => 100, b => 104, p => False, o => False, r => False), (a => 108, b => 112, p => False, o => False, r => False), (a => 116, b => 120, p => False, o => False, r => False), (a => 102, b => 106, p => False, o => False, r => False), (a => 110, b => 114, p => False, o => False, r => False), (a => 118, b => 122, p => False, o => False, r => False), (a => 101, b => 105, p => False, o => False, r => False), (a => 109, b => 113, p => False, o => False, r => False), (a => 117, b => 121, p => False, o => False, r => False), (a => 103, b => 107, p => False, o => False, r => False), (a => 111, b => 115, p => False, o => False, r => False), (a => 119, b => 123, p => False, o => False, r => False), (a => 132, b => 136, p => False, o => False, r => False), (a => 140, b => 144, p => False, o => False, r => False), (a => 148, b => 152, p => False, o => False, r => False), (a => 134, b => 138, p => False, o => False, r => False), (a => 142, b => 146, p => False, o => False, r => False), (a => 150, b => 154, p => False, o => False, r => False), (a => 133, b => 137, p => False, o => False, r => False), (a => 141, b => 145, p => False, o => False, r => False), (a => 149, b => 153, p => False, o => False, r => False), (a => 135, b => 139, p => False, o => False, r => False), (a => 143, b => 147, p => False, o => False, r => False), (a => 151, b => 155, p => False, o => False, r => False), (a => 164, b => 168, p => False, o => False, r => False), (a => 172, b => 176, p => False, o => False, r => False), (a => 180, b => 184, p => False, o => False, r => False), (a => 166, b => 170, p => False, o => False, r => False), (a => 174, b => 178, p => False, o => False, r => False), (a => 182, b => 186, p => False, o => False, r => False), (a => 165, b => 169, p => False, o => False, r => False), (a => 173, b => 177, p => False, o => False, r => False), (a => 181, b => 185, p => False, o => False, r => False), (a => 167, b => 171, p => False, o => False, r => False), (a => 175, b => 179, p => False, o => False, r => False), (a => 183, b => 187, p => False, o => False, r => False), (a => 196, b => 200, p => False, o => False, r => False), (a => 204, b => 208, p => False, o => False, r => False), (a => 212, b => 216, p => False, o => False, r => False), (a => 198, b => 202, p => False, o => False, r => False), (a => 206, b => 210, p => False, o => False, r => False), (a => 214, b => 218, p => False, o => False, r => False), (a => 197, b => 201, p => False, o => False, r => False), (a => 205, b => 209, p => False, o => False, r => False), (a => 213, b => 217, p => False, o => False, r => False), (a => 199, b => 203, p => False, o => False, r => False), (a => 207, b => 211, p => False, o => False, r => False), (a => 215, b => 219, p => False, o => False, r => False), (a => 228, b => 232, p => False, o => False, r => False), (a => 236, b => 240, p => False, o => False, r => False), (a => 244, b => 248, p => False, o => False, r => False), (a => 230, b => 234, p => False, o => False, r => False), (a => 238, b => 242, p => False, o => False, r => False), (a => 246, b => 250, p => False, o => False, r => False), (a => 229, b => 233, p => False, o => False, r => False), (a => 237, b => 241, p => False, o => False, r => False), (a => 245, b => 249, p => False, o => False, r => False), (a => 231, b => 235, p => False, o => False, r => False), (a => 239, b => 243, p => False, o => False, r => False), (a => 247, b => 251, p => False, o => False, r => False), (a => 260, b => 264, p => False, o => False, r => False), (a => 268, b => 272, p => False, o => False, r => False), (a => 276, b => 280, p => False, o => False, r => False), (a => 262, b => 266, p => False, o => False, r => False), (a => 270, b => 274, p => False, o => False, r => False), (a => 278, b => 282, p => False, o => False, r => False), (a => 261, b => 265, p => False, o => False, r => False), (a => 269, b => 273, p => False, o => False, r => False), (a => 277, b => 281, p => False, o => False, r => False), (a => 263, b => 267, p => False, o => False, r => False), (a => 271, b => 275, p => False, o => False, r => False), (a => 279, b => 283, p => False, o => False, r => False), (a => 292, b => 296, p => False, o => False, r => False), (a => 300, b => 304, p => False, o => False, r => False), (a => 308, b => 312, p => False, o => False, r => False), (a => 294, b => 298, p => False, o => False, r => False), (a => 302, b => 306, p => False, o => False, r => False), (a => 310, b => 314, p => False, o => False, r => False), (a => 293, b => 297, p => False, o => False, r => False), (a => 301, b => 305, p => False, o => False, r => False), (a => 309, b => 313, p => False, o => False, r => False), (a => 295, b => 299, p => False, o => False, r => False), (a => 303, b => 307, p => False, o => False, r => False), (a => 311, b => 315, p => False, o => False, r => False), (a => 324, b => 328, p => False, o => False, r => False), (a => 332, b => 336, p => False, o => False, r => False), (a => 340, b => 344, p => False, o => False, r => False), (a => 326, b => 330, p => False, o => False, r => False), (a => 334, b => 338, p => False, o => False, r => False), (a => 342, b => 346, p => False, o => False, r => False), (a => 325, b => 329, p => False, o => False, r => False), (a => 333, b => 337, p => False, o => False, r => False), (a => 341, b => 345, p => False, o => False, r => False), (a => 327, b => 331, p => False, o => False, r => False), (a => 335, b => 339, p => False, o => False, r => False), (a => 343, b => 347, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 28, b => 323, p => True, o => False, r => False), (a => 29, b => 322, p => True, o => False, r => False), (a => 30, b => 321, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 33, b => 318, p => True, o => False, r => False), (a => 34, b => 317, p => True, o => False, r => False), (a => 35, b => 316, p => True, o => False, r => False), (a => 60, b => 291, p => True, o => False, r => False), (a => 61, b => 290, p => True, o => False, r => False), (a => 62, b => 289, p => True, o => False, r => False), (a => 63, b => 288, p => True, o => False, r => False), (a => 64, b => 287, p => True, o => False, r => False), (a => 65, b => 286, p => True, o => False, r => False), (a => 66, b => 285, p => True, o => False, r => False), (a => 67, b => 284, p => True, o => False, r => False), (a => 92, b => 259, p => True, o => False, r => False), (a => 93, b => 258, p => True, o => False, r => False), (a => 94, b => 257, p => True, o => False, r => False), (a => 95, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 98, b => 253, p => True, o => False, r => False), (a => 99, b => 252, p => True, o => False, r => False), (a => 124, b => 227, p => True, o => False, r => False), (a => 125, b => 226, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 129, b => 222, p => True, o => False, r => False), (a => 130, b => 221, p => True, o => False, r => False), (a => 131, b => 220, p => True, o => False, r => False), (a => 156, b => 195, p => True, o => False, r => False), (a => 157, b => 194, p => True, o => False, r => False), (a => 158, b => 193, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 161, b => 190, p => True, o => False, r => False), (a => 162, b => 189, p => True, o => False, r => False), (a => 163, b => 188, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 22, b => 24, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 23, b => 25, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 38, b => 40, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 46, b => 48, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 54, b => 56, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 39, b => 41, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 47, b => 49, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 55, b => 57, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 70, b => 72, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 78, b => 80, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 86, b => 88, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 71, b => 73, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 79, b => 81, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 87, b => 89, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 102, b => 104, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 110, b => 112, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 118, b => 120, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 103, b => 105, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 111, b => 113, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 119, b => 121, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 134, b => 136, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 142, b => 144, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 150, b => 152, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 135, b => 137, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 143, b => 145, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 151, b => 153, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 166, b => 168, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 174, b => 176, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 182, b => 184, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 167, b => 169, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 175, b => 177, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 183, b => 185, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 198, b => 200, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 206, b => 208, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 214, b => 216, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 199, b => 201, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 207, b => 209, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 215, b => 217, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 230, b => 232, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 238, b => 240, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 246, b => 248, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 231, b => 233, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 239, b => 241, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 247, b => 249, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 262, b => 264, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 270, b => 272, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 278, b => 280, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 263, b => 265, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 271, b => 273, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 279, b => 281, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 294, b => 296, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 302, b => 304, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 310, b => 312, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 295, b => 297, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 303, b => 305, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 311, b => 313, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 326, b => 328, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 334, b => 336, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 342, b => 344, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 327, b => 329, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 335, b => 337, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 343, b => 345, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 30, b => 321, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 33, b => 318, p => True, o => False, r => False), (a => 62, b => 289, p => True, o => False, r => False), (a => 63, b => 288, p => True, o => False, r => False), (a => 64, b => 287, p => True, o => False, r => False), (a => 65, b => 286, p => True, o => False, r => False), (a => 94, b => 257, p => True, o => False, r => False), (a => 95, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 129, b => 222, p => True, o => False, r => False), (a => 158, b => 193, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 161, b => 190, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 15, b => 16, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 23, b => 24, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 39, b => 40, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 47, b => 48, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 55, b => 56, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 71, b => 72, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 79, b => 80, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 87, b => 88, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 103, b => 104, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 111, b => 112, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 119, b => 120, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 135, b => 136, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 143, b => 144, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 151, b => 152, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 167, b => 168, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 175, b => 176, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 183, b => 184, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 199, b => 200, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 207, b => 208, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 215, b => 216, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 231, b => 232, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 239, b => 240, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 247, b => 248, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 263, b => 264, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 271, b => 272, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 279, b => 280, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 295, b => 296, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 303, b => 304, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 311, b => 312, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 327, b => 328, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 335, b => 336, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 343, b => 344, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 32, b => 319, p => True, o => False, r => False), (a => 63, b => 288, p => True, o => False, r => False), (a => 64, b => 287, p => True, o => False, r => False), (a => 95, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 223, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False)),
					((a => 16, b => 48, p => False, o => False, r => False), (a => 8, b => 40, p => False, o => False, r => False), (a => 24, b => 56, p => False, o => False, r => False), (a => 4, b => 36, p => False, o => False, r => False), (a => 20, b => 52, p => False, o => False, r => False), (a => 12, b => 44, p => False, o => False, r => False), (a => 28, b => 60, p => False, o => False, r => False), (a => 2, b => 34, p => False, o => False, r => False), (a => 18, b => 50, p => False, o => False, r => False), (a => 10, b => 42, p => False, o => False, r => False), (a => 26, b => 58, p => False, o => False, r => False), (a => 6, b => 38, p => False, o => False, r => False), (a => 22, b => 54, p => False, o => False, r => False), (a => 14, b => 46, p => False, o => False, r => False), (a => 30, b => 62, p => False, o => False, r => False), (a => 1, b => 33, p => False, o => False, r => False), (a => 17, b => 49, p => False, o => False, r => False), (a => 9, b => 41, p => False, o => False, r => False), (a => 25, b => 57, p => False, o => False, r => False), (a => 5, b => 37, p => False, o => False, r => False), (a => 21, b => 53, p => False, o => False, r => False), (a => 13, b => 45, p => False, o => False, r => False), (a => 29, b => 61, p => False, o => False, r => False), (a => 3, b => 35, p => False, o => False, r => False), (a => 19, b => 51, p => False, o => False, r => False), (a => 11, b => 43, p => False, o => False, r => False), (a => 27, b => 59, p => False, o => False, r => False), (a => 7, b => 39, p => False, o => False, r => False), (a => 23, b => 55, p => False, o => False, r => False), (a => 15, b => 47, p => False, o => False, r => False), (a => 80, b => 112, p => False, o => False, r => False), (a => 72, b => 104, p => False, o => False, r => False), (a => 88, b => 120, p => False, o => False, r => False), (a => 68, b => 100, p => False, o => False, r => False), (a => 84, b => 116, p => False, o => False, r => False), (a => 76, b => 108, p => False, o => False, r => False), (a => 92, b => 124, p => False, o => False, r => False), (a => 66, b => 98, p => False, o => False, r => False), (a => 82, b => 114, p => False, o => False, r => False), (a => 74, b => 106, p => False, o => False, r => False), (a => 90, b => 122, p => False, o => False, r => False), (a => 70, b => 102, p => False, o => False, r => False), (a => 86, b => 118, p => False, o => False, r => False), (a => 78, b => 110, p => False, o => False, r => False), (a => 94, b => 126, p => False, o => False, r => False), (a => 65, b => 97, p => False, o => False, r => False), (a => 81, b => 113, p => False, o => False, r => False), (a => 73, b => 105, p => False, o => False, r => False), (a => 89, b => 121, p => False, o => False, r => False), (a => 69, b => 101, p => False, o => False, r => False), (a => 85, b => 117, p => False, o => False, r => False), (a => 77, b => 109, p => False, o => False, r => False), (a => 93, b => 125, p => False, o => False, r => False), (a => 67, b => 99, p => False, o => False, r => False), (a => 83, b => 115, p => False, o => False, r => False), (a => 75, b => 107, p => False, o => False, r => False), (a => 91, b => 123, p => False, o => False, r => False), (a => 71, b => 103, p => False, o => False, r => False), (a => 87, b => 119, p => False, o => False, r => False), (a => 79, b => 111, p => False, o => False, r => False), (a => 144, b => 176, p => False, o => False, r => False), (a => 136, b => 168, p => False, o => False, r => False), (a => 152, b => 184, p => False, o => False, r => False), (a => 132, b => 164, p => False, o => False, r => False), (a => 148, b => 180, p => False, o => False, r => False), (a => 140, b => 172, p => False, o => False, r => False), (a => 156, b => 188, p => False, o => False, r => False), (a => 130, b => 162, p => False, o => False, r => False), (a => 146, b => 178, p => False, o => False, r => False), (a => 138, b => 170, p => False, o => False, r => False), (a => 154, b => 186, p => False, o => False, r => False), (a => 134, b => 166, p => False, o => False, r => False), (a => 150, b => 182, p => False, o => False, r => False), (a => 142, b => 174, p => False, o => False, r => False), (a => 158, b => 190, p => False, o => False, r => False), (a => 129, b => 161, p => False, o => False, r => False), (a => 145, b => 177, p => False, o => False, r => False), (a => 137, b => 169, p => False, o => False, r => False), (a => 153, b => 185, p => False, o => False, r => False), (a => 133, b => 165, p => False, o => False, r => False), (a => 149, b => 181, p => False, o => False, r => False), (a => 141, b => 173, p => False, o => False, r => False), (a => 157, b => 189, p => False, o => False, r => False), (a => 131, b => 163, p => False, o => False, r => False), (a => 147, b => 179, p => False, o => False, r => False), (a => 139, b => 171, p => False, o => False, r => False), (a => 155, b => 187, p => False, o => False, r => False), (a => 135, b => 167, p => False, o => False, r => False), (a => 151, b => 183, p => False, o => False, r => False), (a => 143, b => 175, p => False, o => False, r => False), (a => 208, b => 240, p => False, o => False, r => False), (a => 200, b => 232, p => False, o => False, r => False), (a => 216, b => 248, p => False, o => False, r => False), (a => 196, b => 228, p => False, o => False, r => False), (a => 212, b => 244, p => False, o => False, r => False), (a => 204, b => 236, p => False, o => False, r => False), (a => 220, b => 252, p => False, o => False, r => False), (a => 194, b => 226, p => False, o => False, r => False), (a => 210, b => 242, p => False, o => False, r => False), (a => 202, b => 234, p => False, o => False, r => False), (a => 218, b => 250, p => False, o => False, r => False), (a => 198, b => 230, p => False, o => False, r => False), (a => 214, b => 246, p => False, o => False, r => False), (a => 206, b => 238, p => False, o => False, r => False), (a => 222, b => 254, p => False, o => False, r => False), (a => 193, b => 225, p => False, o => False, r => False), (a => 209, b => 241, p => False, o => False, r => False), (a => 201, b => 233, p => False, o => False, r => False), (a => 217, b => 249, p => False, o => False, r => False), (a => 197, b => 229, p => False, o => False, r => False), (a => 213, b => 245, p => False, o => False, r => False), (a => 205, b => 237, p => False, o => False, r => False), (a => 221, b => 253, p => False, o => False, r => False), (a => 195, b => 227, p => False, o => False, r => False), (a => 211, b => 243, p => False, o => False, r => False), (a => 203, b => 235, p => False, o => False, r => False), (a => 219, b => 251, p => False, o => False, r => False), (a => 199, b => 231, p => False, o => False, r => False), (a => 215, b => 247, p => False, o => False, r => False), (a => 207, b => 239, p => False, o => False, r => False), (a => 272, b => 304, p => False, o => False, r => False), (a => 264, b => 296, p => False, o => False, r => False), (a => 280, b => 312, p => False, o => False, r => False), (a => 260, b => 292, p => False, o => False, r => False), (a => 276, b => 308, p => False, o => False, r => False), (a => 268, b => 300, p => False, o => False, r => False), (a => 284, b => 316, p => False, o => False, r => False), (a => 258, b => 290, p => False, o => False, r => False), (a => 274, b => 306, p => False, o => False, r => False), (a => 266, b => 298, p => False, o => False, r => False), (a => 282, b => 314, p => False, o => False, r => False), (a => 262, b => 294, p => False, o => False, r => False), (a => 278, b => 310, p => False, o => False, r => False), (a => 270, b => 302, p => False, o => False, r => False), (a => 286, b => 318, p => False, o => False, r => False), (a => 257, b => 289, p => False, o => False, r => False), (a => 273, b => 305, p => False, o => False, r => False), (a => 265, b => 297, p => False, o => False, r => False), (a => 281, b => 313, p => False, o => False, r => False), (a => 261, b => 293, p => False, o => False, r => False), (a => 277, b => 309, p => False, o => False, r => False), (a => 269, b => 301, p => False, o => False, r => False), (a => 285, b => 317, p => False, o => False, r => False), (a => 259, b => 291, p => False, o => False, r => False), (a => 275, b => 307, p => False, o => False, r => False), (a => 267, b => 299, p => False, o => False, r => False), (a => 283, b => 315, p => False, o => False, r => False), (a => 263, b => 295, p => False, o => False, r => False), (a => 279, b => 311, p => False, o => False, r => False), (a => 271, b => 303, p => False, o => False, r => False), (a => 328, b => 336, p => False, o => False, r => False), (a => 332, b => 340, p => False, o => False, r => False), (a => 330, b => 338, p => False, o => False, r => False), (a => 334, b => 342, p => False, o => False, r => False), (a => 329, b => 337, p => False, o => False, r => False), (a => 333, b => 341, p => False, o => False, r => False), (a => 331, b => 339, p => False, o => False, r => False), (a => 335, b => 343, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 31, b => 350, p => True, o => False, r => False), (a => 32, b => 349, p => True, o => False, r => False), (a => 63, b => 348, p => True, o => False, r => False), (a => 64, b => 347, p => True, o => False, r => False), (a => 95, b => 346, p => True, o => False, r => False), (a => 96, b => 345, p => True, o => False, r => False), (a => 127, b => 344, p => True, o => False, r => False), (a => 128, b => 327, p => True, o => False, r => False), (a => 159, b => 326, p => True, o => False, r => False), (a => 160, b => 325, p => True, o => False, r => False), (a => 191, b => 324, p => True, o => False, r => False), (a => 192, b => 323, p => True, o => False, r => False), (a => 223, b => 322, p => True, o => False, r => False), (a => 224, b => 321, p => True, o => False, r => False), (a => 255, b => 320, p => True, o => False, r => False), (a => 256, b => 319, p => True, o => False, r => False), (a => 287, b => 288, p => True, o => False, r => False)),
					((a => 16, b => 32, p => False, o => False, r => False), (a => 24, b => 40, p => False, o => False, r => False), (a => 20, b => 36, p => False, o => False, r => False), (a => 28, b => 44, p => False, o => False, r => False), (a => 18, b => 34, p => False, o => False, r => False), (a => 26, b => 42, p => False, o => False, r => False), (a => 22, b => 38, p => False, o => False, r => False), (a => 30, b => 46, p => False, o => False, r => False), (a => 17, b => 33, p => False, o => False, r => False), (a => 25, b => 41, p => False, o => False, r => False), (a => 21, b => 37, p => False, o => False, r => False), (a => 29, b => 45, p => False, o => False, r => False), (a => 19, b => 35, p => False, o => False, r => False), (a => 27, b => 43, p => False, o => False, r => False), (a => 23, b => 39, p => False, o => False, r => False), (a => 31, b => 47, p => False, o => False, r => False), (a => 80, b => 96, p => False, o => False, r => False), (a => 88, b => 104, p => False, o => False, r => False), (a => 84, b => 100, p => False, o => False, r => False), (a => 92, b => 108, p => False, o => False, r => False), (a => 82, b => 98, p => False, o => False, r => False), (a => 90, b => 106, p => False, o => False, r => False), (a => 86, b => 102, p => False, o => False, r => False), (a => 94, b => 110, p => False, o => False, r => False), (a => 81, b => 97, p => False, o => False, r => False), (a => 89, b => 105, p => False, o => False, r => False), (a => 85, b => 101, p => False, o => False, r => False), (a => 93, b => 109, p => False, o => False, r => False), (a => 83, b => 99, p => False, o => False, r => False), (a => 91, b => 107, p => False, o => False, r => False), (a => 87, b => 103, p => False, o => False, r => False), (a => 95, b => 111, p => False, o => False, r => False), (a => 144, b => 160, p => False, o => False, r => False), (a => 152, b => 168, p => False, o => False, r => False), (a => 148, b => 164, p => False, o => False, r => False), (a => 156, b => 172, p => False, o => False, r => False), (a => 146, b => 162, p => False, o => False, r => False), (a => 154, b => 170, p => False, o => False, r => False), (a => 150, b => 166, p => False, o => False, r => False), (a => 158, b => 174, p => False, o => False, r => False), (a => 145, b => 161, p => False, o => False, r => False), (a => 153, b => 169, p => False, o => False, r => False), (a => 149, b => 165, p => False, o => False, r => False), (a => 157, b => 173, p => False, o => False, r => False), (a => 147, b => 163, p => False, o => False, r => False), (a => 155, b => 171, p => False, o => False, r => False), (a => 151, b => 167, p => False, o => False, r => False), (a => 159, b => 175, p => False, o => False, r => False), (a => 208, b => 224, p => False, o => False, r => False), (a => 216, b => 232, p => False, o => False, r => False), (a => 212, b => 228, p => False, o => False, r => False), (a => 220, b => 236, p => False, o => False, r => False), (a => 210, b => 226, p => False, o => False, r => False), (a => 218, b => 234, p => False, o => False, r => False), (a => 214, b => 230, p => False, o => False, r => False), (a => 222, b => 238, p => False, o => False, r => False), (a => 209, b => 225, p => False, o => False, r => False), (a => 217, b => 233, p => False, o => False, r => False), (a => 213, b => 229, p => False, o => False, r => False), (a => 221, b => 237, p => False, o => False, r => False), (a => 211, b => 227, p => False, o => False, r => False), (a => 219, b => 235, p => False, o => False, r => False), (a => 215, b => 231, p => False, o => False, r => False), (a => 223, b => 239, p => False, o => False, r => False), (a => 272, b => 288, p => False, o => False, r => False), (a => 280, b => 296, p => False, o => False, r => False), (a => 276, b => 292, p => False, o => False, r => False), (a => 284, b => 300, p => False, o => False, r => False), (a => 274, b => 290, p => False, o => False, r => False), (a => 282, b => 298, p => False, o => False, r => False), (a => 278, b => 294, p => False, o => False, r => False), (a => 286, b => 302, p => False, o => False, r => False), (a => 273, b => 289, p => False, o => False, r => False), (a => 281, b => 297, p => False, o => False, r => False), (a => 277, b => 293, p => False, o => False, r => False), (a => 285, b => 301, p => False, o => False, r => False), (a => 275, b => 291, p => False, o => False, r => False), (a => 283, b => 299, p => False, o => False, r => False), (a => 279, b => 295, p => False, o => False, r => False), (a => 287, b => 303, p => False, o => False, r => False), (a => 324, b => 328, p => False, o => False, r => False), (a => 332, b => 336, p => False, o => False, r => False), (a => 340, b => 344, p => False, o => False, r => False), (a => 326, b => 330, p => False, o => False, r => False), (a => 334, b => 338, p => False, o => False, r => False), (a => 342, b => 346, p => False, o => False, r => False), (a => 325, b => 329, p => False, o => False, r => False), (a => 333, b => 337, p => False, o => False, r => False), (a => 341, b => 345, p => False, o => False, r => False), (a => 327, b => 331, p => False, o => False, r => False), (a => 335, b => 339, p => False, o => False, r => False), (a => 343, b => 347, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 323, p => True, o => False, r => False), (a => 5, b => 322, p => True, o => False, r => False), (a => 6, b => 321, p => True, o => False, r => False), (a => 7, b => 320, p => True, o => False, r => False), (a => 8, b => 319, p => True, o => False, r => False), (a => 9, b => 318, p => True, o => False, r => False), (a => 10, b => 317, p => True, o => False, r => False), (a => 11, b => 316, p => True, o => False, r => False), (a => 12, b => 315, p => True, o => False, r => False), (a => 13, b => 314, p => True, o => False, r => False), (a => 14, b => 313, p => True, o => False, r => False), (a => 15, b => 312, p => True, o => False, r => False), (a => 48, b => 311, p => True, o => False, r => False), (a => 49, b => 310, p => True, o => False, r => False), (a => 50, b => 309, p => True, o => False, r => False), (a => 51, b => 308, p => True, o => False, r => False), (a => 52, b => 307, p => True, o => False, r => False), (a => 53, b => 306, p => True, o => False, r => False), (a => 54, b => 305, p => True, o => False, r => False), (a => 55, b => 304, p => True, o => False, r => False), (a => 56, b => 271, p => True, o => False, r => False), (a => 57, b => 270, p => True, o => False, r => False), (a => 58, b => 269, p => True, o => False, r => False), (a => 59, b => 268, p => True, o => False, r => False), (a => 60, b => 267, p => True, o => False, r => False), (a => 61, b => 266, p => True, o => False, r => False), (a => 62, b => 265, p => True, o => False, r => False), (a => 63, b => 264, p => True, o => False, r => False), (a => 64, b => 263, p => True, o => False, r => False), (a => 65, b => 262, p => True, o => False, r => False), (a => 66, b => 261, p => True, o => False, r => False), (a => 67, b => 260, p => True, o => False, r => False), (a => 68, b => 259, p => True, o => False, r => False), (a => 69, b => 258, p => True, o => False, r => False), (a => 70, b => 257, p => True, o => False, r => False), (a => 71, b => 256, p => True, o => False, r => False), (a => 72, b => 255, p => True, o => False, r => False), (a => 73, b => 254, p => True, o => False, r => False), (a => 74, b => 253, p => True, o => False, r => False), (a => 75, b => 252, p => True, o => False, r => False), (a => 76, b => 251, p => True, o => False, r => False), (a => 77, b => 250, p => True, o => False, r => False), (a => 78, b => 249, p => True, o => False, r => False), (a => 79, b => 248, p => True, o => False, r => False), (a => 112, b => 247, p => True, o => False, r => False), (a => 113, b => 246, p => True, o => False, r => False), (a => 114, b => 245, p => True, o => False, r => False), (a => 115, b => 244, p => True, o => False, r => False), (a => 116, b => 243, p => True, o => False, r => False), (a => 117, b => 242, p => True, o => False, r => False), (a => 118, b => 241, p => True, o => False, r => False), (a => 119, b => 240, p => True, o => False, r => False), (a => 120, b => 207, p => True, o => False, r => False), (a => 121, b => 206, p => True, o => False, r => False), (a => 122, b => 205, p => True, o => False, r => False), (a => 123, b => 204, p => True, o => False, r => False), (a => 124, b => 203, p => True, o => False, r => False), (a => 125, b => 202, p => True, o => False, r => False), (a => 126, b => 201, p => True, o => False, r => False), (a => 127, b => 200, p => True, o => False, r => False), (a => 128, b => 199, p => True, o => False, r => False), (a => 129, b => 198, p => True, o => False, r => False), (a => 130, b => 197, p => True, o => False, r => False), (a => 131, b => 196, p => True, o => False, r => False), (a => 132, b => 195, p => True, o => False, r => False), (a => 133, b => 194, p => True, o => False, r => False), (a => 134, b => 193, p => True, o => False, r => False), (a => 135, b => 192, p => True, o => False, r => False), (a => 136, b => 191, p => True, o => False, r => False), (a => 137, b => 190, p => True, o => False, r => False), (a => 138, b => 189, p => True, o => False, r => False), (a => 139, b => 188, p => True, o => False, r => False), (a => 140, b => 187, p => True, o => False, r => False), (a => 141, b => 186, p => True, o => False, r => False), (a => 142, b => 185, p => True, o => False, r => False), (a => 143, b => 184, p => True, o => False, r => False), (a => 176, b => 183, p => True, o => False, r => False), (a => 177, b => 182, p => True, o => False, r => False), (a => 178, b => 181, p => True, o => False, r => False), (a => 179, b => 180, p => True, o => False, r => False)),
					((a => 8, b => 16, p => False, o => False, r => False), (a => 24, b => 32, p => False, o => False, r => False), (a => 40, b => 48, p => False, o => False, r => False), (a => 12, b => 20, p => False, o => False, r => False), (a => 28, b => 36, p => False, o => False, r => False), (a => 44, b => 52, p => False, o => False, r => False), (a => 10, b => 18, p => False, o => False, r => False), (a => 26, b => 34, p => False, o => False, r => False), (a => 42, b => 50, p => False, o => False, r => False), (a => 14, b => 22, p => False, o => False, r => False), (a => 30, b => 38, p => False, o => False, r => False), (a => 46, b => 54, p => False, o => False, r => False), (a => 9, b => 17, p => False, o => False, r => False), (a => 25, b => 33, p => False, o => False, r => False), (a => 41, b => 49, p => False, o => False, r => False), (a => 13, b => 21, p => False, o => False, r => False), (a => 29, b => 37, p => False, o => False, r => False), (a => 45, b => 53, p => False, o => False, r => False), (a => 11, b => 19, p => False, o => False, r => False), (a => 27, b => 35, p => False, o => False, r => False), (a => 43, b => 51, p => False, o => False, r => False), (a => 15, b => 23, p => False, o => False, r => False), (a => 31, b => 39, p => False, o => False, r => False), (a => 47, b => 55, p => False, o => False, r => False), (a => 72, b => 80, p => False, o => False, r => False), (a => 88, b => 96, p => False, o => False, r => False), (a => 104, b => 112, p => False, o => False, r => False), (a => 76, b => 84, p => False, o => False, r => False), (a => 92, b => 100, p => False, o => False, r => False), (a => 108, b => 116, p => False, o => False, r => False), (a => 74, b => 82, p => False, o => False, r => False), (a => 90, b => 98, p => False, o => False, r => False), (a => 106, b => 114, p => False, o => False, r => False), (a => 78, b => 86, p => False, o => False, r => False), (a => 94, b => 102, p => False, o => False, r => False), (a => 110, b => 118, p => False, o => False, r => False), (a => 73, b => 81, p => False, o => False, r => False), (a => 89, b => 97, p => False, o => False, r => False), (a => 105, b => 113, p => False, o => False, r => False), (a => 77, b => 85, p => False, o => False, r => False), (a => 93, b => 101, p => False, o => False, r => False), (a => 109, b => 117, p => False, o => False, r => False), (a => 75, b => 83, p => False, o => False, r => False), (a => 91, b => 99, p => False, o => False, r => False), (a => 107, b => 115, p => False, o => False, r => False), (a => 79, b => 87, p => False, o => False, r => False), (a => 95, b => 103, p => False, o => False, r => False), (a => 111, b => 119, p => False, o => False, r => False), (a => 136, b => 144, p => False, o => False, r => False), (a => 152, b => 160, p => False, o => False, r => False), (a => 168, b => 176, p => False, o => False, r => False), (a => 140, b => 148, p => False, o => False, r => False), (a => 156, b => 164, p => False, o => False, r => False), (a => 172, b => 180, p => False, o => False, r => False), (a => 138, b => 146, p => False, o => False, r => False), (a => 154, b => 162, p => False, o => False, r => False), (a => 170, b => 178, p => False, o => False, r => False), (a => 142, b => 150, p => False, o => False, r => False), (a => 158, b => 166, p => False, o => False, r => False), (a => 174, b => 182, p => False, o => False, r => False), (a => 137, b => 145, p => False, o => False, r => False), (a => 153, b => 161, p => False, o => False, r => False), (a => 169, b => 177, p => False, o => False, r => False), (a => 141, b => 149, p => False, o => False, r => False), (a => 157, b => 165, p => False, o => False, r => False), (a => 173, b => 181, p => False, o => False, r => False), (a => 139, b => 147, p => False, o => False, r => False), (a => 155, b => 163, p => False, o => False, r => False), (a => 171, b => 179, p => False, o => False, r => False), (a => 143, b => 151, p => False, o => False, r => False), (a => 159, b => 167, p => False, o => False, r => False), (a => 175, b => 183, p => False, o => False, r => False), (a => 200, b => 208, p => False, o => False, r => False), (a => 216, b => 224, p => False, o => False, r => False), (a => 232, b => 240, p => False, o => False, r => False), (a => 204, b => 212, p => False, o => False, r => False), (a => 220, b => 228, p => False, o => False, r => False), (a => 236, b => 244, p => False, o => False, r => False), (a => 202, b => 210, p => False, o => False, r => False), (a => 218, b => 226, p => False, o => False, r => False), (a => 234, b => 242, p => False, o => False, r => False), (a => 206, b => 214, p => False, o => False, r => False), (a => 222, b => 230, p => False, o => False, r => False), (a => 238, b => 246, p => False, o => False, r => False), (a => 201, b => 209, p => False, o => False, r => False), (a => 217, b => 225, p => False, o => False, r => False), (a => 233, b => 241, p => False, o => False, r => False), (a => 205, b => 213, p => False, o => False, r => False), (a => 221, b => 229, p => False, o => False, r => False), (a => 237, b => 245, p => False, o => False, r => False), (a => 203, b => 211, p => False, o => False, r => False), (a => 219, b => 227, p => False, o => False, r => False), (a => 235, b => 243, p => False, o => False, r => False), (a => 207, b => 215, p => False, o => False, r => False), (a => 223, b => 231, p => False, o => False, r => False), (a => 239, b => 247, p => False, o => False, r => False), (a => 264, b => 272, p => False, o => False, r => False), (a => 280, b => 288, p => False, o => False, r => False), (a => 296, b => 304, p => False, o => False, r => False), (a => 268, b => 276, p => False, o => False, r => False), (a => 284, b => 292, p => False, o => False, r => False), (a => 300, b => 308, p => False, o => False, r => False), (a => 266, b => 274, p => False, o => False, r => False), (a => 282, b => 290, p => False, o => False, r => False), (a => 298, b => 306, p => False, o => False, r => False), (a => 270, b => 278, p => False, o => False, r => False), (a => 286, b => 294, p => False, o => False, r => False), (a => 302, b => 310, p => False, o => False, r => False), (a => 265, b => 273, p => False, o => False, r => False), (a => 281, b => 289, p => False, o => False, r => False), (a => 297, b => 305, p => False, o => False, r => False), (a => 269, b => 277, p => False, o => False, r => False), (a => 285, b => 293, p => False, o => False, r => False), (a => 301, b => 309, p => False, o => False, r => False), (a => 267, b => 275, p => False, o => False, r => False), (a => 283, b => 291, p => False, o => False, r => False), (a => 299, b => 307, p => False, o => False, r => False), (a => 271, b => 279, p => False, o => False, r => False), (a => 287, b => 295, p => False, o => False, r => False), (a => 303, b => 311, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 326, b => 328, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 334, b => 336, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 342, b => 344, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 327, b => 329, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 335, b => 337, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 343, b => 345, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 321, p => True, o => False, r => False), (a => 3, b => 320, p => True, o => False, r => False), (a => 4, b => 319, p => True, o => False, r => False), (a => 5, b => 318, p => True, o => False, r => False), (a => 6, b => 317, p => True, o => False, r => False), (a => 7, b => 316, p => True, o => False, r => False), (a => 56, b => 315, p => True, o => False, r => False), (a => 57, b => 314, p => True, o => False, r => False), (a => 58, b => 313, p => True, o => False, r => False), (a => 59, b => 312, p => True, o => False, r => False), (a => 60, b => 263, p => True, o => False, r => False), (a => 61, b => 262, p => True, o => False, r => False), (a => 62, b => 261, p => True, o => False, r => False), (a => 63, b => 260, p => True, o => False, r => False), (a => 64, b => 259, p => True, o => False, r => False), (a => 65, b => 258, p => True, o => False, r => False), (a => 66, b => 257, p => True, o => False, r => False), (a => 67, b => 256, p => True, o => False, r => False), (a => 68, b => 255, p => True, o => False, r => False), (a => 69, b => 254, p => True, o => False, r => False), (a => 70, b => 253, p => True, o => False, r => False), (a => 71, b => 252, p => True, o => False, r => False), (a => 120, b => 251, p => True, o => False, r => False), (a => 121, b => 250, p => True, o => False, r => False), (a => 122, b => 249, p => True, o => False, r => False), (a => 123, b => 248, p => True, o => False, r => False), (a => 124, b => 199, p => True, o => False, r => False), (a => 125, b => 198, p => True, o => False, r => False), (a => 126, b => 197, p => True, o => False, r => False), (a => 127, b => 196, p => True, o => False, r => False), (a => 128, b => 195, p => True, o => False, r => False), (a => 129, b => 194, p => True, o => False, r => False), (a => 130, b => 193, p => True, o => False, r => False), (a => 131, b => 192, p => True, o => False, r => False), (a => 132, b => 191, p => True, o => False, r => False), (a => 133, b => 190, p => True, o => False, r => False), (a => 134, b => 189, p => True, o => False, r => False), (a => 135, b => 188, p => True, o => False, r => False), (a => 184, b => 187, p => True, o => False, r => False), (a => 185, b => 186, p => True, o => False, r => False)),
					((a => 4, b => 8, p => False, o => False, r => False), (a => 12, b => 16, p => False, o => False, r => False), (a => 20, b => 24, p => False, o => False, r => False), (a => 28, b => 32, p => False, o => False, r => False), (a => 36, b => 40, p => False, o => False, r => False), (a => 44, b => 48, p => False, o => False, r => False), (a => 52, b => 56, p => False, o => False, r => False), (a => 6, b => 10, p => False, o => False, r => False), (a => 14, b => 18, p => False, o => False, r => False), (a => 22, b => 26, p => False, o => False, r => False), (a => 30, b => 34, p => False, o => False, r => False), (a => 38, b => 42, p => False, o => False, r => False), (a => 46, b => 50, p => False, o => False, r => False), (a => 54, b => 58, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 13, b => 17, p => False, o => False, r => False), (a => 21, b => 25, p => False, o => False, r => False), (a => 29, b => 33, p => False, o => False, r => False), (a => 37, b => 41, p => False, o => False, r => False), (a => 45, b => 49, p => False, o => False, r => False), (a => 53, b => 57, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 15, b => 19, p => False, o => False, r => False), (a => 23, b => 27, p => False, o => False, r => False), (a => 31, b => 35, p => False, o => False, r => False), (a => 39, b => 43, p => False, o => False, r => False), (a => 47, b => 51, p => False, o => False, r => False), (a => 55, b => 59, p => False, o => False, r => False), (a => 68, b => 72, p => False, o => False, r => False), (a => 76, b => 80, p => False, o => False, r => False), (a => 84, b => 88, p => False, o => False, r => False), (a => 92, b => 96, p => False, o => False, r => False), (a => 100, b => 104, p => False, o => False, r => False), (a => 108, b => 112, p => False, o => False, r => False), (a => 116, b => 120, p => False, o => False, r => False), (a => 70, b => 74, p => False, o => False, r => False), (a => 78, b => 82, p => False, o => False, r => False), (a => 86, b => 90, p => False, o => False, r => False), (a => 94, b => 98, p => False, o => False, r => False), (a => 102, b => 106, p => False, o => False, r => False), (a => 110, b => 114, p => False, o => False, r => False), (a => 118, b => 122, p => False, o => False, r => False), (a => 69, b => 73, p => False, o => False, r => False), (a => 77, b => 81, p => False, o => False, r => False), (a => 85, b => 89, p => False, o => False, r => False), (a => 93, b => 97, p => False, o => False, r => False), (a => 101, b => 105, p => False, o => False, r => False), (a => 109, b => 113, p => False, o => False, r => False), (a => 117, b => 121, p => False, o => False, r => False), (a => 71, b => 75, p => False, o => False, r => False), (a => 79, b => 83, p => False, o => False, r => False), (a => 87, b => 91, p => False, o => False, r => False), (a => 95, b => 99, p => False, o => False, r => False), (a => 103, b => 107, p => False, o => False, r => False), (a => 111, b => 115, p => False, o => False, r => False), (a => 119, b => 123, p => False, o => False, r => False), (a => 132, b => 136, p => False, o => False, r => False), (a => 140, b => 144, p => False, o => False, r => False), (a => 148, b => 152, p => False, o => False, r => False), (a => 156, b => 160, p => False, o => False, r => False), (a => 164, b => 168, p => False, o => False, r => False), (a => 172, b => 176, p => False, o => False, r => False), (a => 180, b => 184, p => False, o => False, r => False), (a => 134, b => 138, p => False, o => False, r => False), (a => 142, b => 146, p => False, o => False, r => False), (a => 150, b => 154, p => False, o => False, r => False), (a => 158, b => 162, p => False, o => False, r => False), (a => 166, b => 170, p => False, o => False, r => False), (a => 174, b => 178, p => False, o => False, r => False), (a => 182, b => 186, p => False, o => False, r => False), (a => 133, b => 137, p => False, o => False, r => False), (a => 141, b => 145, p => False, o => False, r => False), (a => 149, b => 153, p => False, o => False, r => False), (a => 157, b => 161, p => False, o => False, r => False), (a => 165, b => 169, p => False, o => False, r => False), (a => 173, b => 177, p => False, o => False, r => False), (a => 181, b => 185, p => False, o => False, r => False), (a => 135, b => 139, p => False, o => False, r => False), (a => 143, b => 147, p => False, o => False, r => False), (a => 151, b => 155, p => False, o => False, r => False), (a => 159, b => 163, p => False, o => False, r => False), (a => 167, b => 171, p => False, o => False, r => False), (a => 175, b => 179, p => False, o => False, r => False), (a => 183, b => 187, p => False, o => False, r => False), (a => 196, b => 200, p => False, o => False, r => False), (a => 204, b => 208, p => False, o => False, r => False), (a => 212, b => 216, p => False, o => False, r => False), (a => 220, b => 224, p => False, o => False, r => False), (a => 228, b => 232, p => False, o => False, r => False), (a => 236, b => 240, p => False, o => False, r => False), (a => 244, b => 248, p => False, o => False, r => False), (a => 198, b => 202, p => False, o => False, r => False), (a => 206, b => 210, p => False, o => False, r => False), (a => 214, b => 218, p => False, o => False, r => False), (a => 222, b => 226, p => False, o => False, r => False), (a => 230, b => 234, p => False, o => False, r => False), (a => 238, b => 242, p => False, o => False, r => False), (a => 246, b => 250, p => False, o => False, r => False), (a => 197, b => 201, p => False, o => False, r => False), (a => 205, b => 209, p => False, o => False, r => False), (a => 213, b => 217, p => False, o => False, r => False), (a => 221, b => 225, p => False, o => False, r => False), (a => 229, b => 233, p => False, o => False, r => False), (a => 237, b => 241, p => False, o => False, r => False), (a => 245, b => 249, p => False, o => False, r => False), (a => 199, b => 203, p => False, o => False, r => False), (a => 207, b => 211, p => False, o => False, r => False), (a => 215, b => 219, p => False, o => False, r => False), (a => 223, b => 227, p => False, o => False, r => False), (a => 231, b => 235, p => False, o => False, r => False), (a => 239, b => 243, p => False, o => False, r => False), (a => 247, b => 251, p => False, o => False, r => False), (a => 260, b => 264, p => False, o => False, r => False), (a => 268, b => 272, p => False, o => False, r => False), (a => 276, b => 280, p => False, o => False, r => False), (a => 284, b => 288, p => False, o => False, r => False), (a => 292, b => 296, p => False, o => False, r => False), (a => 300, b => 304, p => False, o => False, r => False), (a => 308, b => 312, p => False, o => False, r => False), (a => 262, b => 266, p => False, o => False, r => False), (a => 270, b => 274, p => False, o => False, r => False), (a => 278, b => 282, p => False, o => False, r => False), (a => 286, b => 290, p => False, o => False, r => False), (a => 294, b => 298, p => False, o => False, r => False), (a => 302, b => 306, p => False, o => False, r => False), (a => 310, b => 314, p => False, o => False, r => False), (a => 261, b => 265, p => False, o => False, r => False), (a => 269, b => 273, p => False, o => False, r => False), (a => 277, b => 281, p => False, o => False, r => False), (a => 285, b => 289, p => False, o => False, r => False), (a => 293, b => 297, p => False, o => False, r => False), (a => 301, b => 305, p => False, o => False, r => False), (a => 309, b => 313, p => False, o => False, r => False), (a => 263, b => 267, p => False, o => False, r => False), (a => 271, b => 275, p => False, o => False, r => False), (a => 279, b => 283, p => False, o => False, r => False), (a => 287, b => 291, p => False, o => False, r => False), (a => 295, b => 299, p => False, o => False, r => False), (a => 303, b => 307, p => False, o => False, r => False), (a => 311, b => 315, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 327, b => 328, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 335, b => 336, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 343, b => 344, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 320, p => True, o => False, r => False), (a => 2, b => 319, p => True, o => False, r => False), (a => 3, b => 318, p => True, o => False, r => False), (a => 60, b => 317, p => True, o => False, r => False), (a => 61, b => 316, p => True, o => False, r => False), (a => 62, b => 259, p => True, o => False, r => False), (a => 63, b => 258, p => True, o => False, r => False), (a => 64, b => 257, p => True, o => False, r => False), (a => 65, b => 256, p => True, o => False, r => False), (a => 66, b => 255, p => True, o => False, r => False), (a => 67, b => 254, p => True, o => False, r => False), (a => 124, b => 253, p => True, o => False, r => False), (a => 125, b => 252, p => True, o => False, r => False), (a => 126, b => 195, p => True, o => False, r => False), (a => 127, b => 194, p => True, o => False, r => False), (a => 128, b => 193, p => True, o => False, r => False), (a => 129, b => 192, p => True, o => False, r => False), (a => 130, b => 191, p => True, o => False, r => False), (a => 131, b => 190, p => True, o => False, r => False), (a => 188, b => 189, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 22, b => 24, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 30, b => 32, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 38, b => 40, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 46, b => 48, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 54, b => 56, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 23, b => 25, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 31, b => 33, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 39, b => 41, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 47, b => 49, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 55, b => 57, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 70, b => 72, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 78, b => 80, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 86, b => 88, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 94, b => 96, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 102, b => 104, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 110, b => 112, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 118, b => 120, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 71, b => 73, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 79, b => 81, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 87, b => 89, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 95, b => 97, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 103, b => 105, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 111, b => 113, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 119, b => 121, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 134, b => 136, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 142, b => 144, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 150, b => 152, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 158, b => 160, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 166, b => 168, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 174, b => 176, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 182, b => 184, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 135, b => 137, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 143, b => 145, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 151, b => 153, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 159, b => 161, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 167, b => 169, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 175, b => 177, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 183, b => 185, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 198, b => 200, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 206, b => 208, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 214, b => 216, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 222, b => 224, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 230, b => 232, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 238, b => 240, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 246, b => 248, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 199, b => 201, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 207, b => 209, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 215, b => 217, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 223, b => 225, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 231, b => 233, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 239, b => 241, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 247, b => 249, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 262, b => 264, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 270, b => 272, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 278, b => 280, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 286, b => 288, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 294, b => 296, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 302, b => 304, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 310, b => 312, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 263, b => 265, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 271, b => 273, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 279, b => 281, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 287, b => 289, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 295, b => 297, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 303, b => 305, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 311, b => 313, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 62, b => 349, p => True, o => False, r => False), (a => 63, b => 348, p => True, o => False, r => False), (a => 64, b => 347, p => True, o => False, r => False), (a => 65, b => 346, p => True, o => False, r => False), (a => 126, b => 345, p => True, o => False, r => False), (a => 127, b => 344, p => True, o => False, r => False), (a => 128, b => 343, p => True, o => False, r => False), (a => 129, b => 342, p => True, o => False, r => False), (a => 190, b => 341, p => True, o => False, r => False), (a => 191, b => 340, p => True, o => False, r => False), (a => 192, b => 339, p => True, o => False, r => False), (a => 193, b => 338, p => True, o => False, r => False), (a => 254, b => 337, p => True, o => False, r => False), (a => 255, b => 336, p => True, o => False, r => False), (a => 256, b => 335, p => True, o => False, r => False), (a => 257, b => 334, p => True, o => False, r => False), (a => 318, b => 333, p => True, o => False, r => False), (a => 319, b => 332, p => True, o => False, r => False), (a => 320, b => 331, p => True, o => False, r => False), (a => 321, b => 330, p => True, o => False, r => False), (a => 322, b => 329, p => True, o => False, r => False), (a => 323, b => 328, p => True, o => False, r => False), (a => 324, b => 327, p => True, o => False, r => False), (a => 325, b => 326, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 15, b => 16, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 23, b => 24, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 31, b => 32, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 39, b => 40, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 47, b => 48, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 55, b => 56, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 71, b => 72, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 79, b => 80, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 87, b => 88, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 95, b => 96, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 103, b => 104, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 111, b => 112, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 119, b => 120, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 135, b => 136, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 143, b => 144, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 151, b => 152, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 159, b => 160, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 167, b => 168, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 175, b => 176, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 183, b => 184, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 199, b => 200, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 207, b => 208, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 215, b => 216, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 223, b => 224, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 231, b => 232, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 239, b => 240, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 247, b => 248, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 263, b => 264, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 271, b => 272, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 279, b => 280, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 287, b => 288, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 295, b => 296, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 303, b => 304, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 311, b => 312, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 63, b => 350, p => True, o => False, r => False), (a => 64, b => 349, p => True, o => False, r => False), (a => 127, b => 348, p => True, o => False, r => False), (a => 128, b => 347, p => True, o => False, r => False), (a => 191, b => 346, p => True, o => False, r => False), (a => 192, b => 345, p => True, o => False, r => False), (a => 255, b => 344, p => True, o => False, r => False), (a => 256, b => 343, p => True, o => False, r => False), (a => 319, b => 342, p => True, o => False, r => False), (a => 320, b => 341, p => True, o => False, r => False), (a => 321, b => 340, p => True, o => False, r => False), (a => 322, b => 339, p => True, o => False, r => False), (a => 323, b => 338, p => True, o => False, r => False), (a => 324, b => 337, p => True, o => False, r => False), (a => 325, b => 336, p => True, o => False, r => False), (a => 326, b => 335, p => True, o => False, r => False), (a => 327, b => 334, p => True, o => False, r => False), (a => 328, b => 333, p => True, o => False, r => False), (a => 329, b => 332, p => True, o => False, r => False), (a => 330, b => 331, p => True, o => False, r => False)),
					((a => 32, b => 96, p => False, o => False, r => False), (a => 16, b => 80, p => False, o => False, r => False), (a => 48, b => 112, p => False, o => False, r => False), (a => 8, b => 72, p => False, o => False, r => False), (a => 40, b => 104, p => False, o => False, r => False), (a => 24, b => 88, p => False, o => False, r => False), (a => 56, b => 120, p => False, o => False, r => False), (a => 4, b => 68, p => False, o => False, r => False), (a => 36, b => 100, p => False, o => False, r => False), (a => 20, b => 84, p => False, o => False, r => False), (a => 52, b => 116, p => False, o => False, r => False), (a => 12, b => 76, p => False, o => False, r => False), (a => 44, b => 108, p => False, o => False, r => False), (a => 28, b => 92, p => False, o => False, r => False), (a => 60, b => 124, p => False, o => False, r => False), (a => 2, b => 66, p => False, o => False, r => False), (a => 34, b => 98, p => False, o => False, r => False), (a => 18, b => 82, p => False, o => False, r => False), (a => 50, b => 114, p => False, o => False, r => False), (a => 10, b => 74, p => False, o => False, r => False), (a => 42, b => 106, p => False, o => False, r => False), (a => 26, b => 90, p => False, o => False, r => False), (a => 58, b => 122, p => False, o => False, r => False), (a => 6, b => 70, p => False, o => False, r => False), (a => 38, b => 102, p => False, o => False, r => False), (a => 22, b => 86, p => False, o => False, r => False), (a => 54, b => 118, p => False, o => False, r => False), (a => 14, b => 78, p => False, o => False, r => False), (a => 46, b => 110, p => False, o => False, r => False), (a => 30, b => 94, p => False, o => False, r => False), (a => 62, b => 126, p => False, o => False, r => False), (a => 1, b => 65, p => False, o => False, r => False), (a => 33, b => 97, p => False, o => False, r => False), (a => 17, b => 81, p => False, o => False, r => False), (a => 49, b => 113, p => False, o => False, r => False), (a => 9, b => 73, p => False, o => False, r => False), (a => 41, b => 105, p => False, o => False, r => False), (a => 25, b => 89, p => False, o => False, r => False), (a => 57, b => 121, p => False, o => False, r => False), (a => 5, b => 69, p => False, o => False, r => False), (a => 37, b => 101, p => False, o => False, r => False), (a => 21, b => 85, p => False, o => False, r => False), (a => 53, b => 117, p => False, o => False, r => False), (a => 13, b => 77, p => False, o => False, r => False), (a => 45, b => 109, p => False, o => False, r => False), (a => 29, b => 93, p => False, o => False, r => False), (a => 61, b => 125, p => False, o => False, r => False), (a => 3, b => 67, p => False, o => False, r => False), (a => 35, b => 99, p => False, o => False, r => False), (a => 19, b => 83, p => False, o => False, r => False), (a => 51, b => 115, p => False, o => False, r => False), (a => 11, b => 75, p => False, o => False, r => False), (a => 43, b => 107, p => False, o => False, r => False), (a => 27, b => 91, p => False, o => False, r => False), (a => 59, b => 123, p => False, o => False, r => False), (a => 7, b => 71, p => False, o => False, r => False), (a => 39, b => 103, p => False, o => False, r => False), (a => 23, b => 87, p => False, o => False, r => False), (a => 55, b => 119, p => False, o => False, r => False), (a => 15, b => 79, p => False, o => False, r => False), (a => 47, b => 111, p => False, o => False, r => False), (a => 31, b => 95, p => False, o => False, r => False), (a => 160, b => 224, p => False, o => False, r => False), (a => 144, b => 208, p => False, o => False, r => False), (a => 176, b => 240, p => False, o => False, r => False), (a => 136, b => 200, p => False, o => False, r => False), (a => 168, b => 232, p => False, o => False, r => False), (a => 152, b => 216, p => False, o => False, r => False), (a => 184, b => 248, p => False, o => False, r => False), (a => 132, b => 196, p => False, o => False, r => False), (a => 164, b => 228, p => False, o => False, r => False), (a => 148, b => 212, p => False, o => False, r => False), (a => 180, b => 244, p => False, o => False, r => False), (a => 140, b => 204, p => False, o => False, r => False), (a => 172, b => 236, p => False, o => False, r => False), (a => 156, b => 220, p => False, o => False, r => False), (a => 188, b => 252, p => False, o => False, r => False), (a => 130, b => 194, p => False, o => False, r => False), (a => 162, b => 226, p => False, o => False, r => False), (a => 146, b => 210, p => False, o => False, r => False), (a => 178, b => 242, p => False, o => False, r => False), (a => 138, b => 202, p => False, o => False, r => False), (a => 170, b => 234, p => False, o => False, r => False), (a => 154, b => 218, p => False, o => False, r => False), (a => 186, b => 250, p => False, o => False, r => False), (a => 134, b => 198, p => False, o => False, r => False), (a => 166, b => 230, p => False, o => False, r => False), (a => 150, b => 214, p => False, o => False, r => False), (a => 182, b => 246, p => False, o => False, r => False), (a => 142, b => 206, p => False, o => False, r => False), (a => 174, b => 238, p => False, o => False, r => False), (a => 158, b => 222, p => False, o => False, r => False), (a => 190, b => 254, p => False, o => False, r => False), (a => 129, b => 193, p => False, o => False, r => False), (a => 161, b => 225, p => False, o => False, r => False), (a => 145, b => 209, p => False, o => False, r => False), (a => 177, b => 241, p => False, o => False, r => False), (a => 137, b => 201, p => False, o => False, r => False), (a => 169, b => 233, p => False, o => False, r => False), (a => 153, b => 217, p => False, o => False, r => False), (a => 185, b => 249, p => False, o => False, r => False), (a => 133, b => 197, p => False, o => False, r => False), (a => 165, b => 229, p => False, o => False, r => False), (a => 149, b => 213, p => False, o => False, r => False), (a => 181, b => 245, p => False, o => False, r => False), (a => 141, b => 205, p => False, o => False, r => False), (a => 173, b => 237, p => False, o => False, r => False), (a => 157, b => 221, p => False, o => False, r => False), (a => 189, b => 253, p => False, o => False, r => False), (a => 131, b => 195, p => False, o => False, r => False), (a => 163, b => 227, p => False, o => False, r => False), (a => 147, b => 211, p => False, o => False, r => False), (a => 179, b => 243, p => False, o => False, r => False), (a => 139, b => 203, p => False, o => False, r => False), (a => 171, b => 235, p => False, o => False, r => False), (a => 155, b => 219, p => False, o => False, r => False), (a => 187, b => 251, p => False, o => False, r => False), (a => 135, b => 199, p => False, o => False, r => False), (a => 167, b => 231, p => False, o => False, r => False), (a => 151, b => 215, p => False, o => False, r => False), (a => 183, b => 247, p => False, o => False, r => False), (a => 143, b => 207, p => False, o => False, r => False), (a => 175, b => 239, p => False, o => False, r => False), (a => 159, b => 223, p => False, o => False, r => False), (a => 288, b => 320, p => False, o => False, r => False), (a => 272, b => 336, p => False, o => False, r => False), (a => 264, b => 328, p => False, o => False, r => False), (a => 280, b => 344, p => False, o => False, r => False), (a => 260, b => 324, p => False, o => False, r => False), (a => 276, b => 340, p => False, o => False, r => False), (a => 268, b => 332, p => False, o => False, r => False), (a => 284, b => 348, p => False, o => False, r => False), (a => 258, b => 322, p => False, o => False, r => False), (a => 274, b => 338, p => False, o => False, r => False), (a => 266, b => 330, p => False, o => False, r => False), (a => 282, b => 346, p => False, o => False, r => False), (a => 262, b => 326, p => False, o => False, r => False), (a => 278, b => 342, p => False, o => False, r => False), (a => 270, b => 334, p => False, o => False, r => False), (a => 286, b => 350, p => False, o => False, r => False), (a => 257, b => 321, p => False, o => False, r => False), (a => 273, b => 337, p => False, o => False, r => False), (a => 265, b => 329, p => False, o => False, r => False), (a => 281, b => 345, p => False, o => False, r => False), (a => 261, b => 325, p => False, o => False, r => False), (a => 277, b => 341, p => False, o => False, r => False), (a => 269, b => 333, p => False, o => False, r => False), (a => 285, b => 349, p => False, o => False, r => False), (a => 259, b => 323, p => False, o => False, r => False), (a => 275, b => 339, p => False, o => False, r => False), (a => 267, b => 331, p => False, o => False, r => False), (a => 283, b => 347, p => False, o => False, r => False), (a => 263, b => 327, p => False, o => False, r => False), (a => 279, b => 343, p => False, o => False, r => False), (a => 271, b => 335, p => False, o => False, r => False), (a => 287, b => 351, p => False, o => False, r => False), (a => 0, b => 319, p => True, o => False, r => False), (a => 63, b => 318, p => True, o => False, r => False), (a => 64, b => 317, p => True, o => False, r => False), (a => 127, b => 316, p => True, o => False, r => False), (a => 128, b => 315, p => True, o => False, r => False), (a => 191, b => 314, p => True, o => False, r => False), (a => 192, b => 313, p => True, o => False, r => False), (a => 255, b => 312, p => True, o => False, r => False), (a => 256, b => 311, p => True, o => False, r => False), (a => 289, b => 310, p => True, o => False, r => False), (a => 290, b => 309, p => True, o => False, r => False), (a => 291, b => 308, p => True, o => False, r => False), (a => 292, b => 307, p => True, o => False, r => False), (a => 293, b => 306, p => True, o => False, r => False), (a => 294, b => 305, p => True, o => False, r => False), (a => 295, b => 304, p => True, o => False, r => False), (a => 296, b => 303, p => True, o => False, r => False), (a => 297, b => 302, p => True, o => False, r => False), (a => 298, b => 301, p => True, o => False, r => False), (a => 299, b => 300, p => True, o => False, r => False)),
					((a => 32, b => 64, p => False, o => False, r => False), (a => 48, b => 80, p => False, o => False, r => False), (a => 40, b => 72, p => False, o => False, r => False), (a => 56, b => 88, p => False, o => False, r => False), (a => 36, b => 68, p => False, o => False, r => False), (a => 52, b => 84, p => False, o => False, r => False), (a => 44, b => 76, p => False, o => False, r => False), (a => 60, b => 92, p => False, o => False, r => False), (a => 34, b => 66, p => False, o => False, r => False), (a => 50, b => 82, p => False, o => False, r => False), (a => 42, b => 74, p => False, o => False, r => False), (a => 58, b => 90, p => False, o => False, r => False), (a => 38, b => 70, p => False, o => False, r => False), (a => 54, b => 86, p => False, o => False, r => False), (a => 46, b => 78, p => False, o => False, r => False), (a => 62, b => 94, p => False, o => False, r => False), (a => 33, b => 65, p => False, o => False, r => False), (a => 49, b => 81, p => False, o => False, r => False), (a => 41, b => 73, p => False, o => False, r => False), (a => 57, b => 89, p => False, o => False, r => False), (a => 37, b => 69, p => False, o => False, r => False), (a => 53, b => 85, p => False, o => False, r => False), (a => 45, b => 77, p => False, o => False, r => False), (a => 61, b => 93, p => False, o => False, r => False), (a => 35, b => 67, p => False, o => False, r => False), (a => 51, b => 83, p => False, o => False, r => False), (a => 43, b => 75, p => False, o => False, r => False), (a => 59, b => 91, p => False, o => False, r => False), (a => 39, b => 71, p => False, o => False, r => False), (a => 55, b => 87, p => False, o => False, r => False), (a => 47, b => 79, p => False, o => False, r => False), (a => 63, b => 95, p => False, o => False, r => False), (a => 160, b => 192, p => False, o => False, r => False), (a => 176, b => 208, p => False, o => False, r => False), (a => 168, b => 200, p => False, o => False, r => False), (a => 184, b => 216, p => False, o => False, r => False), (a => 164, b => 196, p => False, o => False, r => False), (a => 180, b => 212, p => False, o => False, r => False), (a => 172, b => 204, p => False, o => False, r => False), (a => 188, b => 220, p => False, o => False, r => False), (a => 162, b => 194, p => False, o => False, r => False), (a => 178, b => 210, p => False, o => False, r => False), (a => 170, b => 202, p => False, o => False, r => False), (a => 186, b => 218, p => False, o => False, r => False), (a => 166, b => 198, p => False, o => False, r => False), (a => 182, b => 214, p => False, o => False, r => False), (a => 174, b => 206, p => False, o => False, r => False), (a => 190, b => 222, p => False, o => False, r => False), (a => 161, b => 193, p => False, o => False, r => False), (a => 177, b => 209, p => False, o => False, r => False), (a => 169, b => 201, p => False, o => False, r => False), (a => 185, b => 217, p => False, o => False, r => False), (a => 165, b => 197, p => False, o => False, r => False), (a => 181, b => 213, p => False, o => False, r => False), (a => 173, b => 205, p => False, o => False, r => False), (a => 189, b => 221, p => False, o => False, r => False), (a => 163, b => 195, p => False, o => False, r => False), (a => 179, b => 211, p => False, o => False, r => False), (a => 171, b => 203, p => False, o => False, r => False), (a => 187, b => 219, p => False, o => False, r => False), (a => 167, b => 199, p => False, o => False, r => False), (a => 183, b => 215, p => False, o => False, r => False), (a => 175, b => 207, p => False, o => False, r => False), (a => 191, b => 223, p => False, o => False, r => False), (a => 304, b => 336, p => False, o => False, r => False), (a => 272, b => 288, p => False, o => False, r => False), (a => 296, b => 328, p => False, o => False, r => False), (a => 312, b => 344, p => False, o => False, r => False), (a => 292, b => 324, p => False, o => False, r => False), (a => 308, b => 340, p => False, o => False, r => False), (a => 300, b => 332, p => False, o => False, r => False), (a => 316, b => 348, p => False, o => False, r => False), (a => 290, b => 322, p => False, o => False, r => False), (a => 306, b => 338, p => False, o => False, r => False), (a => 298, b => 330, p => False, o => False, r => False), (a => 314, b => 346, p => False, o => False, r => False), (a => 294, b => 326, p => False, o => False, r => False), (a => 310, b => 342, p => False, o => False, r => False), (a => 302, b => 334, p => False, o => False, r => False), (a => 318, b => 350, p => False, o => False, r => False), (a => 289, b => 321, p => False, o => False, r => False), (a => 305, b => 337, p => False, o => False, r => False), (a => 297, b => 329, p => False, o => False, r => False), (a => 313, b => 345, p => False, o => False, r => False), (a => 293, b => 325, p => False, o => False, r => False), (a => 309, b => 341, p => False, o => False, r => False), (a => 301, b => 333, p => False, o => False, r => False), (a => 317, b => 349, p => False, o => False, r => False), (a => 291, b => 323, p => False, o => False, r => False), (a => 307, b => 339, p => False, o => False, r => False), (a => 299, b => 331, p => False, o => False, r => False), (a => 315, b => 347, p => False, o => False, r => False), (a => 295, b => 327, p => False, o => False, r => False), (a => 311, b => 343, p => False, o => False, r => False), (a => 303, b => 335, p => False, o => False, r => False), (a => 319, b => 351, p => False, o => False, r => False), (a => 0, b => 320, p => True, o => False, r => False), (a => 1, b => 287, p => True, o => False, r => False), (a => 2, b => 286, p => True, o => False, r => False), (a => 3, b => 285, p => True, o => False, r => False), (a => 4, b => 284, p => True, o => False, r => False), (a => 5, b => 283, p => True, o => False, r => False), (a => 6, b => 282, p => True, o => False, r => False), (a => 7, b => 281, p => True, o => False, r => False), (a => 8, b => 280, p => True, o => False, r => False), (a => 9, b => 279, p => True, o => False, r => False), (a => 10, b => 278, p => True, o => False, r => False), (a => 11, b => 277, p => True, o => False, r => False), (a => 12, b => 276, p => True, o => False, r => False), (a => 13, b => 275, p => True, o => False, r => False), (a => 14, b => 274, p => True, o => False, r => False), (a => 15, b => 273, p => True, o => False, r => False), (a => 16, b => 271, p => True, o => False, r => False), (a => 17, b => 270, p => True, o => False, r => False), (a => 18, b => 269, p => True, o => False, r => False), (a => 19, b => 268, p => True, o => False, r => False), (a => 20, b => 267, p => True, o => False, r => False), (a => 21, b => 266, p => True, o => False, r => False), (a => 22, b => 265, p => True, o => False, r => False), (a => 23, b => 264, p => True, o => False, r => False), (a => 24, b => 263, p => True, o => False, r => False), (a => 25, b => 262, p => True, o => False, r => False), (a => 26, b => 261, p => True, o => False, r => False), (a => 27, b => 260, p => True, o => False, r => False), (a => 28, b => 259, p => True, o => False, r => False), (a => 29, b => 258, p => True, o => False, r => False), (a => 30, b => 257, p => True, o => False, r => False), (a => 31, b => 256, p => True, o => False, r => False), (a => 96, b => 255, p => True, o => False, r => False), (a => 97, b => 254, p => True, o => False, r => False), (a => 98, b => 253, p => True, o => False, r => False), (a => 99, b => 252, p => True, o => False, r => False), (a => 100, b => 251, p => True, o => False, r => False), (a => 101, b => 250, p => True, o => False, r => False), (a => 102, b => 249, p => True, o => False, r => False), (a => 103, b => 248, p => True, o => False, r => False), (a => 104, b => 247, p => True, o => False, r => False), (a => 105, b => 246, p => True, o => False, r => False), (a => 106, b => 245, p => True, o => False, r => False), (a => 107, b => 244, p => True, o => False, r => False), (a => 108, b => 243, p => True, o => False, r => False), (a => 109, b => 242, p => True, o => False, r => False), (a => 110, b => 241, p => True, o => False, r => False), (a => 111, b => 240, p => True, o => False, r => False), (a => 112, b => 239, p => True, o => False, r => False), (a => 113, b => 238, p => True, o => False, r => False), (a => 114, b => 237, p => True, o => False, r => False), (a => 115, b => 236, p => True, o => False, r => False), (a => 116, b => 235, p => True, o => False, r => False), (a => 117, b => 234, p => True, o => False, r => False), (a => 118, b => 233, p => True, o => False, r => False), (a => 119, b => 232, p => True, o => False, r => False), (a => 120, b => 231, p => True, o => False, r => False), (a => 121, b => 230, p => True, o => False, r => False), (a => 122, b => 229, p => True, o => False, r => False), (a => 123, b => 228, p => True, o => False, r => False), (a => 124, b => 227, p => True, o => False, r => False), (a => 125, b => 226, p => True, o => False, r => False), (a => 126, b => 225, p => True, o => False, r => False), (a => 127, b => 224, p => True, o => False, r => False), (a => 128, b => 159, p => True, o => False, r => False), (a => 129, b => 158, p => True, o => False, r => False), (a => 130, b => 157, p => True, o => False, r => False), (a => 131, b => 156, p => True, o => False, r => False), (a => 132, b => 155, p => True, o => False, r => False), (a => 133, b => 154, p => True, o => False, r => False), (a => 134, b => 153, p => True, o => False, r => False), (a => 135, b => 152, p => True, o => False, r => False), (a => 136, b => 151, p => True, o => False, r => False), (a => 137, b => 150, p => True, o => False, r => False), (a => 138, b => 149, p => True, o => False, r => False), (a => 139, b => 148, p => True, o => False, r => False), (a => 140, b => 147, p => True, o => False, r => False), (a => 141, b => 146, p => True, o => False, r => False), (a => 142, b => 145, p => True, o => False, r => False), (a => 143, b => 144, p => True, o => False, r => False)),
					((a => 16, b => 32, p => False, o => False, r => False), (a => 48, b => 64, p => False, o => False, r => False), (a => 80, b => 96, p => False, o => False, r => False), (a => 24, b => 40, p => False, o => False, r => False), (a => 56, b => 72, p => False, o => False, r => False), (a => 88, b => 104, p => False, o => False, r => False), (a => 20, b => 36, p => False, o => False, r => False), (a => 52, b => 68, p => False, o => False, r => False), (a => 84, b => 100, p => False, o => False, r => False), (a => 28, b => 44, p => False, o => False, r => False), (a => 60, b => 76, p => False, o => False, r => False), (a => 92, b => 108, p => False, o => False, r => False), (a => 18, b => 34, p => False, o => False, r => False), (a => 50, b => 66, p => False, o => False, r => False), (a => 82, b => 98, p => False, o => False, r => False), (a => 26, b => 42, p => False, o => False, r => False), (a => 58, b => 74, p => False, o => False, r => False), (a => 90, b => 106, p => False, o => False, r => False), (a => 22, b => 38, p => False, o => False, r => False), (a => 54, b => 70, p => False, o => False, r => False), (a => 86, b => 102, p => False, o => False, r => False), (a => 30, b => 46, p => False, o => False, r => False), (a => 62, b => 78, p => False, o => False, r => False), (a => 94, b => 110, p => False, o => False, r => False), (a => 17, b => 33, p => False, o => False, r => False), (a => 49, b => 65, p => False, o => False, r => False), (a => 81, b => 97, p => False, o => False, r => False), (a => 25, b => 41, p => False, o => False, r => False), (a => 57, b => 73, p => False, o => False, r => False), (a => 89, b => 105, p => False, o => False, r => False), (a => 21, b => 37, p => False, o => False, r => False), (a => 53, b => 69, p => False, o => False, r => False), (a => 85, b => 101, p => False, o => False, r => False), (a => 29, b => 45, p => False, o => False, r => False), (a => 61, b => 77, p => False, o => False, r => False), (a => 93, b => 109, p => False, o => False, r => False), (a => 19, b => 35, p => False, o => False, r => False), (a => 51, b => 67, p => False, o => False, r => False), (a => 83, b => 99, p => False, o => False, r => False), (a => 27, b => 43, p => False, o => False, r => False), (a => 59, b => 75, p => False, o => False, r => False), (a => 91, b => 107, p => False, o => False, r => False), (a => 23, b => 39, p => False, o => False, r => False), (a => 55, b => 71, p => False, o => False, r => False), (a => 87, b => 103, p => False, o => False, r => False), (a => 31, b => 47, p => False, o => False, r => False), (a => 63, b => 79, p => False, o => False, r => False), (a => 95, b => 111, p => False, o => False, r => False), (a => 144, b => 160, p => False, o => False, r => False), (a => 176, b => 192, p => False, o => False, r => False), (a => 208, b => 224, p => False, o => False, r => False), (a => 152, b => 168, p => False, o => False, r => False), (a => 184, b => 200, p => False, o => False, r => False), (a => 216, b => 232, p => False, o => False, r => False), (a => 148, b => 164, p => False, o => False, r => False), (a => 180, b => 196, p => False, o => False, r => False), (a => 212, b => 228, p => False, o => False, r => False), (a => 156, b => 172, p => False, o => False, r => False), (a => 188, b => 204, p => False, o => False, r => False), (a => 220, b => 236, p => False, o => False, r => False), (a => 146, b => 162, p => False, o => False, r => False), (a => 178, b => 194, p => False, o => False, r => False), (a => 210, b => 226, p => False, o => False, r => False), (a => 154, b => 170, p => False, o => False, r => False), (a => 186, b => 202, p => False, o => False, r => False), (a => 218, b => 234, p => False, o => False, r => False), (a => 150, b => 166, p => False, o => False, r => False), (a => 182, b => 198, p => False, o => False, r => False), (a => 214, b => 230, p => False, o => False, r => False), (a => 158, b => 174, p => False, o => False, r => False), (a => 190, b => 206, p => False, o => False, r => False), (a => 222, b => 238, p => False, o => False, r => False), (a => 145, b => 161, p => False, o => False, r => False), (a => 177, b => 193, p => False, o => False, r => False), (a => 209, b => 225, p => False, o => False, r => False), (a => 153, b => 169, p => False, o => False, r => False), (a => 185, b => 201, p => False, o => False, r => False), (a => 217, b => 233, p => False, o => False, r => False), (a => 149, b => 165, p => False, o => False, r => False), (a => 181, b => 197, p => False, o => False, r => False), (a => 213, b => 229, p => False, o => False, r => False), (a => 157, b => 173, p => False, o => False, r => False), (a => 189, b => 205, p => False, o => False, r => False), (a => 221, b => 237, p => False, o => False, r => False), (a => 147, b => 163, p => False, o => False, r => False), (a => 179, b => 195, p => False, o => False, r => False), (a => 211, b => 227, p => False, o => False, r => False), (a => 155, b => 171, p => False, o => False, r => False), (a => 187, b => 203, p => False, o => False, r => False), (a => 219, b => 235, p => False, o => False, r => False), (a => 151, b => 167, p => False, o => False, r => False), (a => 183, b => 199, p => False, o => False, r => False), (a => 215, b => 231, p => False, o => False, r => False), (a => 159, b => 175, p => False, o => False, r => False), (a => 191, b => 207, p => False, o => False, r => False), (a => 223, b => 239, p => False, o => False, r => False), (a => 304, b => 320, p => False, o => False, r => False), (a => 280, b => 296, p => False, o => False, r => False), (a => 312, b => 328, p => False, o => False, r => False), (a => 264, b => 272, p => False, o => False, r => False), (a => 276, b => 292, p => False, o => False, r => False), (a => 308, b => 324, p => False, o => False, r => False), (a => 284, b => 300, p => False, o => False, r => False), (a => 316, b => 332, p => False, o => False, r => False), (a => 274, b => 290, p => False, o => False, r => False), (a => 306, b => 322, p => False, o => False, r => False), (a => 282, b => 298, p => False, o => False, r => False), (a => 314, b => 330, p => False, o => False, r => False), (a => 278, b => 294, p => False, o => False, r => False), (a => 310, b => 326, p => False, o => False, r => False), (a => 286, b => 302, p => False, o => False, r => False), (a => 318, b => 334, p => False, o => False, r => False), (a => 273, b => 289, p => False, o => False, r => False), (a => 305, b => 321, p => False, o => False, r => False), (a => 281, b => 297, p => False, o => False, r => False), (a => 313, b => 329, p => False, o => False, r => False), (a => 277, b => 293, p => False, o => False, r => False), (a => 309, b => 325, p => False, o => False, r => False), (a => 285, b => 301, p => False, o => False, r => False), (a => 317, b => 333, p => False, o => False, r => False), (a => 275, b => 291, p => False, o => False, r => False), (a => 307, b => 323, p => False, o => False, r => False), (a => 283, b => 299, p => False, o => False, r => False), (a => 315, b => 331, p => False, o => False, r => False), (a => 279, b => 295, p => False, o => False, r => False), (a => 311, b => 327, p => False, o => False, r => False), (a => 287, b => 303, p => False, o => False, r => False), (a => 319, b => 335, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 8, b => 343, p => True, o => False, r => False), (a => 9, b => 342, p => True, o => False, r => False), (a => 10, b => 341, p => True, o => False, r => False), (a => 11, b => 340, p => True, o => False, r => False), (a => 12, b => 339, p => True, o => False, r => False), (a => 13, b => 338, p => True, o => False, r => False), (a => 14, b => 337, p => True, o => False, r => False), (a => 15, b => 336, p => True, o => False, r => False), (a => 112, b => 288, p => True, o => False, r => False), (a => 113, b => 271, p => True, o => False, r => False), (a => 114, b => 270, p => True, o => False, r => False), (a => 115, b => 269, p => True, o => False, r => False), (a => 116, b => 268, p => True, o => False, r => False), (a => 117, b => 267, p => True, o => False, r => False), (a => 118, b => 266, p => True, o => False, r => False), (a => 119, b => 265, p => True, o => False, r => False), (a => 120, b => 263, p => True, o => False, r => False), (a => 121, b => 262, p => True, o => False, r => False), (a => 122, b => 261, p => True, o => False, r => False), (a => 123, b => 260, p => True, o => False, r => False), (a => 124, b => 259, p => True, o => False, r => False), (a => 125, b => 258, p => True, o => False, r => False), (a => 126, b => 257, p => True, o => False, r => False), (a => 127, b => 256, p => True, o => False, r => False), (a => 128, b => 255, p => True, o => False, r => False), (a => 129, b => 254, p => True, o => False, r => False), (a => 130, b => 253, p => True, o => False, r => False), (a => 131, b => 252, p => True, o => False, r => False), (a => 132, b => 251, p => True, o => False, r => False), (a => 133, b => 250, p => True, o => False, r => False), (a => 134, b => 249, p => True, o => False, r => False), (a => 135, b => 248, p => True, o => False, r => False), (a => 136, b => 247, p => True, o => False, r => False), (a => 137, b => 246, p => True, o => False, r => False), (a => 138, b => 245, p => True, o => False, r => False), (a => 139, b => 244, p => True, o => False, r => False), (a => 140, b => 243, p => True, o => False, r => False), (a => 141, b => 242, p => True, o => False, r => False), (a => 142, b => 241, p => True, o => False, r => False), (a => 143, b => 240, p => True, o => False, r => False)),
					((a => 8, b => 16, p => False, o => False, r => False), (a => 24, b => 32, p => False, o => False, r => False), (a => 40, b => 48, p => False, o => False, r => False), (a => 56, b => 64, p => False, o => False, r => False), (a => 72, b => 80, p => False, o => False, r => False), (a => 88, b => 96, p => False, o => False, r => False), (a => 104, b => 112, p => False, o => False, r => False), (a => 12, b => 20, p => False, o => False, r => False), (a => 28, b => 36, p => False, o => False, r => False), (a => 44, b => 52, p => False, o => False, r => False), (a => 60, b => 68, p => False, o => False, r => False), (a => 76, b => 84, p => False, o => False, r => False), (a => 92, b => 100, p => False, o => False, r => False), (a => 108, b => 116, p => False, o => False, r => False), (a => 10, b => 18, p => False, o => False, r => False), (a => 26, b => 34, p => False, o => False, r => False), (a => 42, b => 50, p => False, o => False, r => False), (a => 58, b => 66, p => False, o => False, r => False), (a => 74, b => 82, p => False, o => False, r => False), (a => 90, b => 98, p => False, o => False, r => False), (a => 106, b => 114, p => False, o => False, r => False), (a => 14, b => 22, p => False, o => False, r => False), (a => 30, b => 38, p => False, o => False, r => False), (a => 46, b => 54, p => False, o => False, r => False), (a => 62, b => 70, p => False, o => False, r => False), (a => 78, b => 86, p => False, o => False, r => False), (a => 94, b => 102, p => False, o => False, r => False), (a => 110, b => 118, p => False, o => False, r => False), (a => 9, b => 17, p => False, o => False, r => False), (a => 25, b => 33, p => False, o => False, r => False), (a => 41, b => 49, p => False, o => False, r => False), (a => 57, b => 65, p => False, o => False, r => False), (a => 73, b => 81, p => False, o => False, r => False), (a => 89, b => 97, p => False, o => False, r => False), (a => 105, b => 113, p => False, o => False, r => False), (a => 13, b => 21, p => False, o => False, r => False), (a => 29, b => 37, p => False, o => False, r => False), (a => 45, b => 53, p => False, o => False, r => False), (a => 61, b => 69, p => False, o => False, r => False), (a => 77, b => 85, p => False, o => False, r => False), (a => 93, b => 101, p => False, o => False, r => False), (a => 109, b => 117, p => False, o => False, r => False), (a => 11, b => 19, p => False, o => False, r => False), (a => 27, b => 35, p => False, o => False, r => False), (a => 43, b => 51, p => False, o => False, r => False), (a => 59, b => 67, p => False, o => False, r => False), (a => 75, b => 83, p => False, o => False, r => False), (a => 91, b => 99, p => False, o => False, r => False), (a => 107, b => 115, p => False, o => False, r => False), (a => 15, b => 23, p => False, o => False, r => False), (a => 31, b => 39, p => False, o => False, r => False), (a => 47, b => 55, p => False, o => False, r => False), (a => 63, b => 71, p => False, o => False, r => False), (a => 79, b => 87, p => False, o => False, r => False), (a => 95, b => 103, p => False, o => False, r => False), (a => 111, b => 119, p => False, o => False, r => False), (a => 136, b => 144, p => False, o => False, r => False), (a => 152, b => 160, p => False, o => False, r => False), (a => 168, b => 176, p => False, o => False, r => False), (a => 184, b => 192, p => False, o => False, r => False), (a => 200, b => 208, p => False, o => False, r => False), (a => 216, b => 224, p => False, o => False, r => False), (a => 232, b => 240, p => False, o => False, r => False), (a => 140, b => 148, p => False, o => False, r => False), (a => 156, b => 164, p => False, o => False, r => False), (a => 172, b => 180, p => False, o => False, r => False), (a => 188, b => 196, p => False, o => False, r => False), (a => 204, b => 212, p => False, o => False, r => False), (a => 220, b => 228, p => False, o => False, r => False), (a => 236, b => 244, p => False, o => False, r => False), (a => 138, b => 146, p => False, o => False, r => False), (a => 154, b => 162, p => False, o => False, r => False), (a => 170, b => 178, p => False, o => False, r => False), (a => 186, b => 194, p => False, o => False, r => False), (a => 202, b => 210, p => False, o => False, r => False), (a => 218, b => 226, p => False, o => False, r => False), (a => 234, b => 242, p => False, o => False, r => False), (a => 142, b => 150, p => False, o => False, r => False), (a => 158, b => 166, p => False, o => False, r => False), (a => 174, b => 182, p => False, o => False, r => False), (a => 190, b => 198, p => False, o => False, r => False), (a => 206, b => 214, p => False, o => False, r => False), (a => 222, b => 230, p => False, o => False, r => False), (a => 238, b => 246, p => False, o => False, r => False), (a => 137, b => 145, p => False, o => False, r => False), (a => 153, b => 161, p => False, o => False, r => False), (a => 169, b => 177, p => False, o => False, r => False), (a => 185, b => 193, p => False, o => False, r => False), (a => 201, b => 209, p => False, o => False, r => False), (a => 217, b => 225, p => False, o => False, r => False), (a => 233, b => 241, p => False, o => False, r => False), (a => 141, b => 149, p => False, o => False, r => False), (a => 157, b => 165, p => False, o => False, r => False), (a => 173, b => 181, p => False, o => False, r => False), (a => 189, b => 197, p => False, o => False, r => False), (a => 205, b => 213, p => False, o => False, r => False), (a => 221, b => 229, p => False, o => False, r => False), (a => 237, b => 245, p => False, o => False, r => False), (a => 139, b => 147, p => False, o => False, r => False), (a => 155, b => 163, p => False, o => False, r => False), (a => 171, b => 179, p => False, o => False, r => False), (a => 187, b => 195, p => False, o => False, r => False), (a => 203, b => 211, p => False, o => False, r => False), (a => 219, b => 227, p => False, o => False, r => False), (a => 235, b => 243, p => False, o => False, r => False), (a => 143, b => 151, p => False, o => False, r => False), (a => 159, b => 167, p => False, o => False, r => False), (a => 175, b => 183, p => False, o => False, r => False), (a => 191, b => 199, p => False, o => False, r => False), (a => 207, b => 215, p => False, o => False, r => False), (a => 223, b => 231, p => False, o => False, r => False), (a => 239, b => 247, p => False, o => False, r => False), (a => 280, b => 288, p => False, o => False, r => False), (a => 296, b => 304, p => False, o => False, r => False), (a => 312, b => 320, p => False, o => False, r => False), (a => 328, b => 336, p => False, o => False, r => False), (a => 268, b => 276, p => False, o => False, r => False), (a => 284, b => 292, p => False, o => False, r => False), (a => 300, b => 308, p => False, o => False, r => False), (a => 316, b => 324, p => False, o => False, r => False), (a => 332, b => 340, p => False, o => False, r => False), (a => 260, b => 264, p => False, o => False, r => False), (a => 266, b => 274, p => False, o => False, r => False), (a => 282, b => 290, p => False, o => False, r => False), (a => 298, b => 306, p => False, o => False, r => False), (a => 314, b => 322, p => False, o => False, r => False), (a => 330, b => 338, p => False, o => False, r => False), (a => 270, b => 278, p => False, o => False, r => False), (a => 286, b => 294, p => False, o => False, r => False), (a => 302, b => 310, p => False, o => False, r => False), (a => 318, b => 326, p => False, o => False, r => False), (a => 334, b => 342, p => False, o => False, r => False), (a => 265, b => 273, p => False, o => False, r => False), (a => 281, b => 289, p => False, o => False, r => False), (a => 297, b => 305, p => False, o => False, r => False), (a => 313, b => 321, p => False, o => False, r => False), (a => 329, b => 337, p => False, o => False, r => False), (a => 269, b => 277, p => False, o => False, r => False), (a => 285, b => 293, p => False, o => False, r => False), (a => 301, b => 309, p => False, o => False, r => False), (a => 317, b => 325, p => False, o => False, r => False), (a => 333, b => 341, p => False, o => False, r => False), (a => 267, b => 275, p => False, o => False, r => False), (a => 283, b => 291, p => False, o => False, r => False), (a => 299, b => 307, p => False, o => False, r => False), (a => 315, b => 323, p => False, o => False, r => False), (a => 331, b => 339, p => False, o => False, r => False), (a => 271, b => 279, p => False, o => False, r => False), (a => 287, b => 295, p => False, o => False, r => False), (a => 303, b => 311, p => False, o => False, r => False), (a => 319, b => 327, p => False, o => False, r => False), (a => 335, b => 343, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 120, b => 272, p => True, o => False, r => False), (a => 121, b => 263, p => True, o => False, r => False), (a => 122, b => 262, p => True, o => False, r => False), (a => 123, b => 261, p => True, o => False, r => False), (a => 124, b => 259, p => True, o => False, r => False), (a => 125, b => 258, p => True, o => False, r => False), (a => 126, b => 257, p => True, o => False, r => False), (a => 127, b => 256, p => True, o => False, r => False), (a => 128, b => 255, p => True, o => False, r => False), (a => 129, b => 254, p => True, o => False, r => False), (a => 130, b => 253, p => True, o => False, r => False), (a => 131, b => 252, p => True, o => False, r => False), (a => 132, b => 251, p => True, o => False, r => False), (a => 133, b => 250, p => True, o => False, r => False), (a => 134, b => 249, p => True, o => False, r => False), (a => 135, b => 248, p => True, o => False, r => False)),
					((a => 4, b => 8, p => False, o => False, r => False), (a => 12, b => 16, p => False, o => False, r => False), (a => 20, b => 24, p => False, o => False, r => False), (a => 28, b => 32, p => False, o => False, r => False), (a => 36, b => 40, p => False, o => False, r => False), (a => 44, b => 48, p => False, o => False, r => False), (a => 52, b => 56, p => False, o => False, r => False), (a => 60, b => 64, p => False, o => False, r => False), (a => 68, b => 72, p => False, o => False, r => False), (a => 76, b => 80, p => False, o => False, r => False), (a => 84, b => 88, p => False, o => False, r => False), (a => 92, b => 96, p => False, o => False, r => False), (a => 100, b => 104, p => False, o => False, r => False), (a => 108, b => 112, p => False, o => False, r => False), (a => 116, b => 120, p => False, o => False, r => False), (a => 6, b => 10, p => False, o => False, r => False), (a => 14, b => 18, p => False, o => False, r => False), (a => 22, b => 26, p => False, o => False, r => False), (a => 30, b => 34, p => False, o => False, r => False), (a => 38, b => 42, p => False, o => False, r => False), (a => 46, b => 50, p => False, o => False, r => False), (a => 54, b => 58, p => False, o => False, r => False), (a => 62, b => 66, p => False, o => False, r => False), (a => 70, b => 74, p => False, o => False, r => False), (a => 78, b => 82, p => False, o => False, r => False), (a => 86, b => 90, p => False, o => False, r => False), (a => 94, b => 98, p => False, o => False, r => False), (a => 102, b => 106, p => False, o => False, r => False), (a => 110, b => 114, p => False, o => False, r => False), (a => 118, b => 122, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 13, b => 17, p => False, o => False, r => False), (a => 21, b => 25, p => False, o => False, r => False), (a => 29, b => 33, p => False, o => False, r => False), (a => 37, b => 41, p => False, o => False, r => False), (a => 45, b => 49, p => False, o => False, r => False), (a => 53, b => 57, p => False, o => False, r => False), (a => 61, b => 65, p => False, o => False, r => False), (a => 69, b => 73, p => False, o => False, r => False), (a => 77, b => 81, p => False, o => False, r => False), (a => 85, b => 89, p => False, o => False, r => False), (a => 93, b => 97, p => False, o => False, r => False), (a => 101, b => 105, p => False, o => False, r => False), (a => 109, b => 113, p => False, o => False, r => False), (a => 117, b => 121, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 15, b => 19, p => False, o => False, r => False), (a => 23, b => 27, p => False, o => False, r => False), (a => 31, b => 35, p => False, o => False, r => False), (a => 39, b => 43, p => False, o => False, r => False), (a => 47, b => 51, p => False, o => False, r => False), (a => 55, b => 59, p => False, o => False, r => False), (a => 63, b => 67, p => False, o => False, r => False), (a => 71, b => 75, p => False, o => False, r => False), (a => 79, b => 83, p => False, o => False, r => False), (a => 87, b => 91, p => False, o => False, r => False), (a => 95, b => 99, p => False, o => False, r => False), (a => 103, b => 107, p => False, o => False, r => False), (a => 111, b => 115, p => False, o => False, r => False), (a => 119, b => 123, p => False, o => False, r => False), (a => 132, b => 136, p => False, o => False, r => False), (a => 140, b => 144, p => False, o => False, r => False), (a => 148, b => 152, p => False, o => False, r => False), (a => 156, b => 160, p => False, o => False, r => False), (a => 164, b => 168, p => False, o => False, r => False), (a => 172, b => 176, p => False, o => False, r => False), (a => 180, b => 184, p => False, o => False, r => False), (a => 188, b => 192, p => False, o => False, r => False), (a => 196, b => 200, p => False, o => False, r => False), (a => 204, b => 208, p => False, o => False, r => False), (a => 212, b => 216, p => False, o => False, r => False), (a => 220, b => 224, p => False, o => False, r => False), (a => 228, b => 232, p => False, o => False, r => False), (a => 236, b => 240, p => False, o => False, r => False), (a => 244, b => 248, p => False, o => False, r => False), (a => 134, b => 138, p => False, o => False, r => False), (a => 142, b => 146, p => False, o => False, r => False), (a => 150, b => 154, p => False, o => False, r => False), (a => 158, b => 162, p => False, o => False, r => False), (a => 166, b => 170, p => False, o => False, r => False), (a => 174, b => 178, p => False, o => False, r => False), (a => 182, b => 186, p => False, o => False, r => False), (a => 190, b => 194, p => False, o => False, r => False), (a => 198, b => 202, p => False, o => False, r => False), (a => 206, b => 210, p => False, o => False, r => False), (a => 214, b => 218, p => False, o => False, r => False), (a => 222, b => 226, p => False, o => False, r => False), (a => 230, b => 234, p => False, o => False, r => False), (a => 238, b => 242, p => False, o => False, r => False), (a => 246, b => 250, p => False, o => False, r => False), (a => 133, b => 137, p => False, o => False, r => False), (a => 141, b => 145, p => False, o => False, r => False), (a => 149, b => 153, p => False, o => False, r => False), (a => 157, b => 161, p => False, o => False, r => False), (a => 165, b => 169, p => False, o => False, r => False), (a => 173, b => 177, p => False, o => False, r => False), (a => 181, b => 185, p => False, o => False, r => False), (a => 189, b => 193, p => False, o => False, r => False), (a => 197, b => 201, p => False, o => False, r => False), (a => 205, b => 209, p => False, o => False, r => False), (a => 213, b => 217, p => False, o => False, r => False), (a => 221, b => 225, p => False, o => False, r => False), (a => 229, b => 233, p => False, o => False, r => False), (a => 237, b => 241, p => False, o => False, r => False), (a => 245, b => 249, p => False, o => False, r => False), (a => 135, b => 139, p => False, o => False, r => False), (a => 143, b => 147, p => False, o => False, r => False), (a => 151, b => 155, p => False, o => False, r => False), (a => 159, b => 163, p => False, o => False, r => False), (a => 167, b => 171, p => False, o => False, r => False), (a => 175, b => 179, p => False, o => False, r => False), (a => 183, b => 187, p => False, o => False, r => False), (a => 191, b => 195, p => False, o => False, r => False), (a => 199, b => 203, p => False, o => False, r => False), (a => 207, b => 211, p => False, o => False, r => False), (a => 215, b => 219, p => False, o => False, r => False), (a => 223, b => 227, p => False, o => False, r => False), (a => 231, b => 235, p => False, o => False, r => False), (a => 239, b => 243, p => False, o => False, r => False), (a => 247, b => 251, p => False, o => False, r => False), (a => 268, b => 272, p => False, o => False, r => False), (a => 276, b => 280, p => False, o => False, r => False), (a => 284, b => 288, p => False, o => False, r => False), (a => 292, b => 296, p => False, o => False, r => False), (a => 300, b => 304, p => False, o => False, r => False), (a => 308, b => 312, p => False, o => False, r => False), (a => 316, b => 320, p => False, o => False, r => False), (a => 324, b => 328, p => False, o => False, r => False), (a => 332, b => 336, p => False, o => False, r => False), (a => 340, b => 344, p => False, o => False, r => False), (a => 262, b => 266, p => False, o => False, r => False), (a => 270, b => 274, p => False, o => False, r => False), (a => 278, b => 282, p => False, o => False, r => False), (a => 286, b => 290, p => False, o => False, r => False), (a => 294, b => 298, p => False, o => False, r => False), (a => 302, b => 306, p => False, o => False, r => False), (a => 310, b => 314, p => False, o => False, r => False), (a => 318, b => 322, p => False, o => False, r => False), (a => 326, b => 330, p => False, o => False, r => False), (a => 334, b => 338, p => False, o => False, r => False), (a => 342, b => 346, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 261, b => 265, p => False, o => False, r => False), (a => 269, b => 273, p => False, o => False, r => False), (a => 277, b => 281, p => False, o => False, r => False), (a => 285, b => 289, p => False, o => False, r => False), (a => 293, b => 297, p => False, o => False, r => False), (a => 301, b => 305, p => False, o => False, r => False), (a => 309, b => 313, p => False, o => False, r => False), (a => 317, b => 321, p => False, o => False, r => False), (a => 325, b => 329, p => False, o => False, r => False), (a => 333, b => 337, p => False, o => False, r => False), (a => 341, b => 345, p => False, o => False, r => False), (a => 263, b => 267, p => False, o => False, r => False), (a => 271, b => 275, p => False, o => False, r => False), (a => 279, b => 283, p => False, o => False, r => False), (a => 287, b => 291, p => False, o => False, r => False), (a => 295, b => 299, p => False, o => False, r => False), (a => 303, b => 307, p => False, o => False, r => False), (a => 311, b => 315, p => False, o => False, r => False), (a => 319, b => 323, p => False, o => False, r => False), (a => 327, b => 331, p => False, o => False, r => False), (a => 335, b => 339, p => False, o => False, r => False), (a => 343, b => 347, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 124, b => 264, p => True, o => False, r => False), (a => 125, b => 259, p => True, o => False, r => False), (a => 126, b => 257, p => True, o => False, r => False), (a => 127, b => 256, p => True, o => False, r => False), (a => 128, b => 255, p => True, o => False, r => False), (a => 129, b => 254, p => True, o => False, r => False), (a => 130, b => 253, p => True, o => False, r => False), (a => 131, b => 252, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 22, b => 24, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 30, b => 32, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 38, b => 40, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 46, b => 48, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 54, b => 56, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 62, b => 64, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 70, b => 72, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 78, b => 80, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 86, b => 88, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 94, b => 96, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 102, b => 104, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 110, b => 112, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 118, b => 120, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 23, b => 25, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 31, b => 33, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 39, b => 41, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 47, b => 49, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 55, b => 57, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 63, b => 65, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 71, b => 73, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 79, b => 81, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 87, b => 89, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 95, b => 97, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 103, b => 105, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 111, b => 113, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 119, b => 121, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 134, b => 136, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 142, b => 144, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 150, b => 152, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 158, b => 160, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 166, b => 168, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 174, b => 176, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 182, b => 184, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 190, b => 192, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 198, b => 200, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 206, b => 208, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 214, b => 216, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 222, b => 224, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 230, b => 232, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 238, b => 240, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 246, b => 248, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 135, b => 137, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 143, b => 145, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 151, b => 153, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 159, b => 161, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 167, b => 169, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 175, b => 177, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 183, b => 185, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 191, b => 193, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 199, b => 201, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 207, b => 209, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 215, b => 217, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 223, b => 225, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 231, b => 233, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 239, b => 241, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 247, b => 249, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 262, b => 264, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 270, b => 272, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 278, b => 280, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 286, b => 288, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 294, b => 296, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 302, b => 304, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 310, b => 312, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 318, b => 320, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 326, b => 328, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 334, b => 336, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 342, b => 344, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 263, b => 265, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 271, b => 273, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 279, b => 281, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 287, b => 289, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 295, b => 297, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 303, b => 305, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 311, b => 313, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 319, b => 321, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 327, b => 329, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 335, b => 337, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 343, b => 345, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 126, b => 260, p => True, o => False, r => False), (a => 127, b => 256, p => True, o => False, r => False), (a => 128, b => 255, p => True, o => False, r => False), (a => 129, b => 254, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 15, b => 16, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 23, b => 24, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 31, b => 32, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 39, b => 40, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 47, b => 48, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 55, b => 56, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 63, b => 64, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 71, b => 72, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 79, b => 80, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 87, b => 88, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 95, b => 96, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 103, b => 104, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 111, b => 112, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 119, b => 120, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 135, b => 136, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 143, b => 144, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 151, b => 152, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 159, b => 160, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 167, b => 168, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 175, b => 176, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 183, b => 184, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 191, b => 192, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 199, b => 200, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 207, b => 208, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 215, b => 216, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 223, b => 224, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 231, b => 232, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 239, b => 240, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 247, b => 248, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 263, b => 264, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 271, b => 272, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 279, b => 280, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 287, b => 288, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 295, b => 296, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 303, b => 304, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 311, b => 312, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 319, b => 320, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 327, b => 328, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 335, b => 336, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 343, b => 344, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 127, b => 258, p => True, o => False, r => False), (a => 128, b => 257, p => True, o => False, r => False), (a => 255, b => 256, p => True, o => False, r => False)),
					((a => 64, b => 192, p => False, o => False, r => False), (a => 32, b => 160, p => False, o => False, r => False), (a => 96, b => 224, p => False, o => False, r => False), (a => 16, b => 144, p => False, o => False, r => False), (a => 80, b => 208, p => False, o => False, r => False), (a => 48, b => 176, p => False, o => False, r => False), (a => 112, b => 240, p => False, o => False, r => False), (a => 8, b => 136, p => False, o => False, r => False), (a => 72, b => 200, p => False, o => False, r => False), (a => 40, b => 168, p => False, o => False, r => False), (a => 104, b => 232, p => False, o => False, r => False), (a => 24, b => 152, p => False, o => False, r => False), (a => 88, b => 216, p => False, o => False, r => False), (a => 56, b => 184, p => False, o => False, r => False), (a => 120, b => 248, p => False, o => False, r => False), (a => 4, b => 132, p => False, o => False, r => False), (a => 68, b => 196, p => False, o => False, r => False), (a => 36, b => 164, p => False, o => False, r => False), (a => 100, b => 228, p => False, o => False, r => False), (a => 20, b => 148, p => False, o => False, r => False), (a => 84, b => 212, p => False, o => False, r => False), (a => 52, b => 180, p => False, o => False, r => False), (a => 116, b => 244, p => False, o => False, r => False), (a => 12, b => 140, p => False, o => False, r => False), (a => 76, b => 204, p => False, o => False, r => False), (a => 44, b => 172, p => False, o => False, r => False), (a => 108, b => 236, p => False, o => False, r => False), (a => 28, b => 156, p => False, o => False, r => False), (a => 92, b => 220, p => False, o => False, r => False), (a => 60, b => 188, p => False, o => False, r => False), (a => 124, b => 252, p => False, o => False, r => False), (a => 2, b => 130, p => False, o => False, r => False), (a => 66, b => 194, p => False, o => False, r => False), (a => 34, b => 162, p => False, o => False, r => False), (a => 98, b => 226, p => False, o => False, r => False), (a => 18, b => 146, p => False, o => False, r => False), (a => 82, b => 210, p => False, o => False, r => False), (a => 50, b => 178, p => False, o => False, r => False), (a => 114, b => 242, p => False, o => False, r => False), (a => 10, b => 138, p => False, o => False, r => False), (a => 74, b => 202, p => False, o => False, r => False), (a => 42, b => 170, p => False, o => False, r => False), (a => 106, b => 234, p => False, o => False, r => False), (a => 26, b => 154, p => False, o => False, r => False), (a => 90, b => 218, p => False, o => False, r => False), (a => 58, b => 186, p => False, o => False, r => False), (a => 122, b => 250, p => False, o => False, r => False), (a => 6, b => 134, p => False, o => False, r => False), (a => 70, b => 198, p => False, o => False, r => False), (a => 38, b => 166, p => False, o => False, r => False), (a => 102, b => 230, p => False, o => False, r => False), (a => 22, b => 150, p => False, o => False, r => False), (a => 86, b => 214, p => False, o => False, r => False), (a => 54, b => 182, p => False, o => False, r => False), (a => 118, b => 246, p => False, o => False, r => False), (a => 14, b => 142, p => False, o => False, r => False), (a => 78, b => 206, p => False, o => False, r => False), (a => 46, b => 174, p => False, o => False, r => False), (a => 110, b => 238, p => False, o => False, r => False), (a => 30, b => 158, p => False, o => False, r => False), (a => 94, b => 222, p => False, o => False, r => False), (a => 62, b => 190, p => False, o => False, r => False), (a => 126, b => 254, p => False, o => False, r => False), (a => 1, b => 129, p => False, o => False, r => False), (a => 65, b => 193, p => False, o => False, r => False), (a => 33, b => 161, p => False, o => False, r => False), (a => 97, b => 225, p => False, o => False, r => False), (a => 17, b => 145, p => False, o => False, r => False), (a => 81, b => 209, p => False, o => False, r => False), (a => 49, b => 177, p => False, o => False, r => False), (a => 113, b => 241, p => False, o => False, r => False), (a => 9, b => 137, p => False, o => False, r => False), (a => 73, b => 201, p => False, o => False, r => False), (a => 41, b => 169, p => False, o => False, r => False), (a => 105, b => 233, p => False, o => False, r => False), (a => 25, b => 153, p => False, o => False, r => False), (a => 89, b => 217, p => False, o => False, r => False), (a => 57, b => 185, p => False, o => False, r => False), (a => 121, b => 249, p => False, o => False, r => False), (a => 5, b => 133, p => False, o => False, r => False), (a => 69, b => 197, p => False, o => False, r => False), (a => 37, b => 165, p => False, o => False, r => False), (a => 101, b => 229, p => False, o => False, r => False), (a => 21, b => 149, p => False, o => False, r => False), (a => 85, b => 213, p => False, o => False, r => False), (a => 53, b => 181, p => False, o => False, r => False), (a => 117, b => 245, p => False, o => False, r => False), (a => 13, b => 141, p => False, o => False, r => False), (a => 77, b => 205, p => False, o => False, r => False), (a => 45, b => 173, p => False, o => False, r => False), (a => 109, b => 237, p => False, o => False, r => False), (a => 29, b => 157, p => False, o => False, r => False), (a => 93, b => 221, p => False, o => False, r => False), (a => 61, b => 189, p => False, o => False, r => False), (a => 125, b => 253, p => False, o => False, r => False), (a => 3, b => 131, p => False, o => False, r => False), (a => 67, b => 195, p => False, o => False, r => False), (a => 35, b => 163, p => False, o => False, r => False), (a => 99, b => 227, p => False, o => False, r => False), (a => 19, b => 147, p => False, o => False, r => False), (a => 83, b => 211, p => False, o => False, r => False), (a => 51, b => 179, p => False, o => False, r => False), (a => 115, b => 243, p => False, o => False, r => False), (a => 11, b => 139, p => False, o => False, r => False), (a => 75, b => 203, p => False, o => False, r => False), (a => 43, b => 171, p => False, o => False, r => False), (a => 107, b => 235, p => False, o => False, r => False), (a => 27, b => 155, p => False, o => False, r => False), (a => 91, b => 219, p => False, o => False, r => False), (a => 59, b => 187, p => False, o => False, r => False), (a => 123, b => 251, p => False, o => False, r => False), (a => 7, b => 135, p => False, o => False, r => False), (a => 71, b => 199, p => False, o => False, r => False), (a => 39, b => 167, p => False, o => False, r => False), (a => 103, b => 231, p => False, o => False, r => False), (a => 23, b => 151, p => False, o => False, r => False), (a => 87, b => 215, p => False, o => False, r => False), (a => 55, b => 183, p => False, o => False, r => False), (a => 119, b => 247, p => False, o => False, r => False), (a => 15, b => 143, p => False, o => False, r => False), (a => 79, b => 207, p => False, o => False, r => False), (a => 47, b => 175, p => False, o => False, r => False), (a => 111, b => 239, p => False, o => False, r => False), (a => 31, b => 159, p => False, o => False, r => False), (a => 95, b => 223, p => False, o => False, r => False), (a => 63, b => 191, p => False, o => False, r => False), (a => 288, b => 320, p => False, o => False, r => False), (a => 304, b => 336, p => False, o => False, r => False), (a => 296, b => 328, p => False, o => False, r => False), (a => 312, b => 344, p => False, o => False, r => False), (a => 292, b => 324, p => False, o => False, r => False), (a => 308, b => 340, p => False, o => False, r => False), (a => 300, b => 332, p => False, o => False, r => False), (a => 316, b => 348, p => False, o => False, r => False), (a => 290, b => 322, p => False, o => False, r => False), (a => 306, b => 338, p => False, o => False, r => False), (a => 298, b => 330, p => False, o => False, r => False), (a => 314, b => 346, p => False, o => False, r => False), (a => 294, b => 326, p => False, o => False, r => False), (a => 310, b => 342, p => False, o => False, r => False), (a => 302, b => 334, p => False, o => False, r => False), (a => 318, b => 350, p => False, o => False, r => False), (a => 289, b => 321, p => False, o => False, r => False), (a => 305, b => 337, p => False, o => False, r => False), (a => 297, b => 329, p => False, o => False, r => False), (a => 313, b => 345, p => False, o => False, r => False), (a => 293, b => 325, p => False, o => False, r => False), (a => 309, b => 341, p => False, o => False, r => False), (a => 301, b => 333, p => False, o => False, r => False), (a => 317, b => 349, p => False, o => False, r => False), (a => 291, b => 323, p => False, o => False, r => False), (a => 307, b => 339, p => False, o => False, r => False), (a => 299, b => 331, p => False, o => False, r => False), (a => 315, b => 347, p => False, o => False, r => False), (a => 295, b => 327, p => False, o => False, r => False), (a => 311, b => 343, p => False, o => False, r => False), (a => 303, b => 335, p => False, o => False, r => False), (a => 319, b => 351, p => False, o => False, r => False), (a => 0, b => 287, p => True, o => False, r => False), (a => 127, b => 286, p => True, o => False, r => False), (a => 128, b => 285, p => True, o => False, r => False), (a => 255, b => 284, p => True, o => False, r => False), (a => 256, b => 283, p => True, o => False, r => False), (a => 257, b => 282, p => True, o => False, r => False), (a => 258, b => 281, p => True, o => False, r => False), (a => 259, b => 280, p => True, o => False, r => False), (a => 260, b => 279, p => True, o => False, r => False), (a => 261, b => 278, p => True, o => False, r => False), (a => 262, b => 277, p => True, o => False, r => False), (a => 263, b => 276, p => True, o => False, r => False), (a => 264, b => 275, p => True, o => False, r => False), (a => 265, b => 274, p => True, o => False, r => False), (a => 266, b => 273, p => True, o => False, r => False), (a => 267, b => 272, p => True, o => False, r => False), (a => 268, b => 271, p => True, o => False, r => False), (a => 269, b => 270, p => True, o => False, r => False)),
					((a => 64, b => 128, p => False, o => False, r => False), (a => 96, b => 160, p => False, o => False, r => False), (a => 80, b => 144, p => False, o => False, r => False), (a => 112, b => 176, p => False, o => False, r => False), (a => 72, b => 136, p => False, o => False, r => False), (a => 104, b => 168, p => False, o => False, r => False), (a => 88, b => 152, p => False, o => False, r => False), (a => 120, b => 184, p => False, o => False, r => False), (a => 68, b => 132, p => False, o => False, r => False), (a => 100, b => 164, p => False, o => False, r => False), (a => 84, b => 148, p => False, o => False, r => False), (a => 116, b => 180, p => False, o => False, r => False), (a => 76, b => 140, p => False, o => False, r => False), (a => 108, b => 172, p => False, o => False, r => False), (a => 92, b => 156, p => False, o => False, r => False), (a => 124, b => 188, p => False, o => False, r => False), (a => 66, b => 130, p => False, o => False, r => False), (a => 98, b => 162, p => False, o => False, r => False), (a => 82, b => 146, p => False, o => False, r => False), (a => 114, b => 178, p => False, o => False, r => False), (a => 74, b => 138, p => False, o => False, r => False), (a => 106, b => 170, p => False, o => False, r => False), (a => 90, b => 154, p => False, o => False, r => False), (a => 122, b => 186, p => False, o => False, r => False), (a => 70, b => 134, p => False, o => False, r => False), (a => 102, b => 166, p => False, o => False, r => False), (a => 86, b => 150, p => False, o => False, r => False), (a => 118, b => 182, p => False, o => False, r => False), (a => 78, b => 142, p => False, o => False, r => False), (a => 110, b => 174, p => False, o => False, r => False), (a => 94, b => 158, p => False, o => False, r => False), (a => 126, b => 190, p => False, o => False, r => False), (a => 65, b => 129, p => False, o => False, r => False), (a => 97, b => 161, p => False, o => False, r => False), (a => 81, b => 145, p => False, o => False, r => False), (a => 113, b => 177, p => False, o => False, r => False), (a => 73, b => 137, p => False, o => False, r => False), (a => 105, b => 169, p => False, o => False, r => False), (a => 89, b => 153, p => False, o => False, r => False), (a => 121, b => 185, p => False, o => False, r => False), (a => 69, b => 133, p => False, o => False, r => False), (a => 101, b => 165, p => False, o => False, r => False), (a => 85, b => 149, p => False, o => False, r => False), (a => 117, b => 181, p => False, o => False, r => False), (a => 77, b => 141, p => False, o => False, r => False), (a => 109, b => 173, p => False, o => False, r => False), (a => 93, b => 157, p => False, o => False, r => False), (a => 125, b => 189, p => False, o => False, r => False), (a => 67, b => 131, p => False, o => False, r => False), (a => 99, b => 163, p => False, o => False, r => False), (a => 83, b => 147, p => False, o => False, r => False), (a => 115, b => 179, p => False, o => False, r => False), (a => 75, b => 139, p => False, o => False, r => False), (a => 107, b => 171, p => False, o => False, r => False), (a => 91, b => 155, p => False, o => False, r => False), (a => 123, b => 187, p => False, o => False, r => False), (a => 71, b => 135, p => False, o => False, r => False), (a => 103, b => 167, p => False, o => False, r => False), (a => 87, b => 151, p => False, o => False, r => False), (a => 119, b => 183, p => False, o => False, r => False), (a => 79, b => 143, p => False, o => False, r => False), (a => 111, b => 175, p => False, o => False, r => False), (a => 95, b => 159, p => False, o => False, r => False), (a => 127, b => 191, p => False, o => False, r => False), (a => 272, b => 288, p => False, o => False, r => False), (a => 304, b => 320, p => False, o => False, r => False), (a => 280, b => 296, p => False, o => False, r => False), (a => 312, b => 328, p => False, o => False, r => False), (a => 276, b => 292, p => False, o => False, r => False), (a => 308, b => 324, p => False, o => False, r => False), (a => 284, b => 300, p => False, o => False, r => False), (a => 316, b => 332, p => False, o => False, r => False), (a => 274, b => 290, p => False, o => False, r => False), (a => 306, b => 322, p => False, o => False, r => False), (a => 282, b => 298, p => False, o => False, r => False), (a => 314, b => 330, p => False, o => False, r => False), (a => 278, b => 294, p => False, o => False, r => False), (a => 310, b => 326, p => False, o => False, r => False), (a => 286, b => 302, p => False, o => False, r => False), (a => 318, b => 334, p => False, o => False, r => False), (a => 273, b => 289, p => False, o => False, r => False), (a => 305, b => 321, p => False, o => False, r => False), (a => 281, b => 297, p => False, o => False, r => False), (a => 313, b => 329, p => False, o => False, r => False), (a => 277, b => 293, p => False, o => False, r => False), (a => 309, b => 325, p => False, o => False, r => False), (a => 285, b => 301, p => False, o => False, r => False), (a => 317, b => 333, p => False, o => False, r => False), (a => 275, b => 291, p => False, o => False, r => False), (a => 307, b => 323, p => False, o => False, r => False), (a => 283, b => 299, p => False, o => False, r => False), (a => 315, b => 331, p => False, o => False, r => False), (a => 279, b => 295, p => False, o => False, r => False), (a => 311, b => 327, p => False, o => False, r => False), (a => 287, b => 303, p => False, o => False, r => False), (a => 319, b => 335, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 8, b => 343, p => True, o => False, r => False), (a => 9, b => 342, p => True, o => False, r => False), (a => 10, b => 341, p => True, o => False, r => False), (a => 11, b => 340, p => True, o => False, r => False), (a => 12, b => 339, p => True, o => False, r => False), (a => 13, b => 338, p => True, o => False, r => False), (a => 14, b => 337, p => True, o => False, r => False), (a => 15, b => 336, p => True, o => False, r => False), (a => 16, b => 271, p => True, o => False, r => False), (a => 17, b => 270, p => True, o => False, r => False), (a => 18, b => 269, p => True, o => False, r => False), (a => 19, b => 268, p => True, o => False, r => False), (a => 20, b => 267, p => True, o => False, r => False), (a => 21, b => 266, p => True, o => False, r => False), (a => 22, b => 265, p => True, o => False, r => False), (a => 23, b => 264, p => True, o => False, r => False), (a => 24, b => 263, p => True, o => False, r => False), (a => 25, b => 262, p => True, o => False, r => False), (a => 26, b => 261, p => True, o => False, r => False), (a => 27, b => 260, p => True, o => False, r => False), (a => 28, b => 259, p => True, o => False, r => False), (a => 29, b => 258, p => True, o => False, r => False), (a => 30, b => 257, p => True, o => False, r => False), (a => 31, b => 256, p => True, o => False, r => False), (a => 32, b => 255, p => True, o => False, r => False), (a => 33, b => 254, p => True, o => False, r => False), (a => 34, b => 253, p => True, o => False, r => False), (a => 35, b => 252, p => True, o => False, r => False), (a => 36, b => 251, p => True, o => False, r => False), (a => 37, b => 250, p => True, o => False, r => False), (a => 38, b => 249, p => True, o => False, r => False), (a => 39, b => 248, p => True, o => False, r => False), (a => 40, b => 247, p => True, o => False, r => False), (a => 41, b => 246, p => True, o => False, r => False), (a => 42, b => 245, p => True, o => False, r => False), (a => 43, b => 244, p => True, o => False, r => False), (a => 44, b => 243, p => True, o => False, r => False), (a => 45, b => 242, p => True, o => False, r => False), (a => 46, b => 241, p => True, o => False, r => False), (a => 47, b => 240, p => True, o => False, r => False), (a => 48, b => 239, p => True, o => False, r => False), (a => 49, b => 238, p => True, o => False, r => False), (a => 50, b => 237, p => True, o => False, r => False), (a => 51, b => 236, p => True, o => False, r => False), (a => 52, b => 235, p => True, o => False, r => False), (a => 53, b => 234, p => True, o => False, r => False), (a => 54, b => 233, p => True, o => False, r => False), (a => 55, b => 232, p => True, o => False, r => False), (a => 56, b => 231, p => True, o => False, r => False), (a => 57, b => 230, p => True, o => False, r => False), (a => 58, b => 229, p => True, o => False, r => False), (a => 59, b => 228, p => True, o => False, r => False), (a => 60, b => 227, p => True, o => False, r => False), (a => 61, b => 226, p => True, o => False, r => False), (a => 62, b => 225, p => True, o => False, r => False), (a => 63, b => 224, p => True, o => False, r => False), (a => 192, b => 223, p => True, o => False, r => False), (a => 193, b => 222, p => True, o => False, r => False), (a => 194, b => 221, p => True, o => False, r => False), (a => 195, b => 220, p => True, o => False, r => False), (a => 196, b => 219, p => True, o => False, r => False), (a => 197, b => 218, p => True, o => False, r => False), (a => 198, b => 217, p => True, o => False, r => False), (a => 199, b => 216, p => True, o => False, r => False), (a => 200, b => 215, p => True, o => False, r => False), (a => 201, b => 214, p => True, o => False, r => False), (a => 202, b => 213, p => True, o => False, r => False), (a => 203, b => 212, p => True, o => False, r => False), (a => 204, b => 211, p => True, o => False, r => False), (a => 205, b => 210, p => True, o => False, r => False), (a => 206, b => 209, p => True, o => False, r => False), (a => 207, b => 208, p => True, o => False, r => False)),
					((a => 32, b => 64, p => False, o => False, r => False), (a => 96, b => 128, p => False, o => False, r => False), (a => 160, b => 192, p => False, o => False, r => False), (a => 48, b => 80, p => False, o => False, r => False), (a => 112, b => 144, p => False, o => False, r => False), (a => 176, b => 208, p => False, o => False, r => False), (a => 40, b => 72, p => False, o => False, r => False), (a => 104, b => 136, p => False, o => False, r => False), (a => 168, b => 200, p => False, o => False, r => False), (a => 56, b => 88, p => False, o => False, r => False), (a => 120, b => 152, p => False, o => False, r => False), (a => 184, b => 216, p => False, o => False, r => False), (a => 36, b => 68, p => False, o => False, r => False), (a => 100, b => 132, p => False, o => False, r => False), (a => 164, b => 196, p => False, o => False, r => False), (a => 52, b => 84, p => False, o => False, r => False), (a => 116, b => 148, p => False, o => False, r => False), (a => 180, b => 212, p => False, o => False, r => False), (a => 44, b => 76, p => False, o => False, r => False), (a => 108, b => 140, p => False, o => False, r => False), (a => 172, b => 204, p => False, o => False, r => False), (a => 60, b => 92, p => False, o => False, r => False), (a => 124, b => 156, p => False, o => False, r => False), (a => 188, b => 220, p => False, o => False, r => False), (a => 34, b => 66, p => False, o => False, r => False), (a => 98, b => 130, p => False, o => False, r => False), (a => 162, b => 194, p => False, o => False, r => False), (a => 50, b => 82, p => False, o => False, r => False), (a => 114, b => 146, p => False, o => False, r => False), (a => 178, b => 210, p => False, o => False, r => False), (a => 42, b => 74, p => False, o => False, r => False), (a => 106, b => 138, p => False, o => False, r => False), (a => 170, b => 202, p => False, o => False, r => False), (a => 58, b => 90, p => False, o => False, r => False), (a => 122, b => 154, p => False, o => False, r => False), (a => 186, b => 218, p => False, o => False, r => False), (a => 38, b => 70, p => False, o => False, r => False), (a => 102, b => 134, p => False, o => False, r => False), (a => 166, b => 198, p => False, o => False, r => False), (a => 54, b => 86, p => False, o => False, r => False), (a => 118, b => 150, p => False, o => False, r => False), (a => 182, b => 214, p => False, o => False, r => False), (a => 46, b => 78, p => False, o => False, r => False), (a => 110, b => 142, p => False, o => False, r => False), (a => 174, b => 206, p => False, o => False, r => False), (a => 62, b => 94, p => False, o => False, r => False), (a => 126, b => 158, p => False, o => False, r => False), (a => 190, b => 222, p => False, o => False, r => False), (a => 33, b => 65, p => False, o => False, r => False), (a => 97, b => 129, p => False, o => False, r => False), (a => 161, b => 193, p => False, o => False, r => False), (a => 49, b => 81, p => False, o => False, r => False), (a => 113, b => 145, p => False, o => False, r => False), (a => 177, b => 209, p => False, o => False, r => False), (a => 41, b => 73, p => False, o => False, r => False), (a => 105, b => 137, p => False, o => False, r => False), (a => 169, b => 201, p => False, o => False, r => False), (a => 57, b => 89, p => False, o => False, r => False), (a => 121, b => 153, p => False, o => False, r => False), (a => 185, b => 217, p => False, o => False, r => False), (a => 37, b => 69, p => False, o => False, r => False), (a => 101, b => 133, p => False, o => False, r => False), (a => 165, b => 197, p => False, o => False, r => False), (a => 53, b => 85, p => False, o => False, r => False), (a => 117, b => 149, p => False, o => False, r => False), (a => 181, b => 213, p => False, o => False, r => False), (a => 45, b => 77, p => False, o => False, r => False), (a => 109, b => 141, p => False, o => False, r => False), (a => 173, b => 205, p => False, o => False, r => False), (a => 61, b => 93, p => False, o => False, r => False), (a => 125, b => 157, p => False, o => False, r => False), (a => 189, b => 221, p => False, o => False, r => False), (a => 35, b => 67, p => False, o => False, r => False), (a => 99, b => 131, p => False, o => False, r => False), (a => 163, b => 195, p => False, o => False, r => False), (a => 51, b => 83, p => False, o => False, r => False), (a => 115, b => 147, p => False, o => False, r => False), (a => 179, b => 211, p => False, o => False, r => False), (a => 43, b => 75, p => False, o => False, r => False), (a => 107, b => 139, p => False, o => False, r => False), (a => 171, b => 203, p => False, o => False, r => False), (a => 59, b => 91, p => False, o => False, r => False), (a => 123, b => 155, p => False, o => False, r => False), (a => 187, b => 219, p => False, o => False, r => False), (a => 39, b => 71, p => False, o => False, r => False), (a => 103, b => 135, p => False, o => False, r => False), (a => 167, b => 199, p => False, o => False, r => False), (a => 55, b => 87, p => False, o => False, r => False), (a => 119, b => 151, p => False, o => False, r => False), (a => 183, b => 215, p => False, o => False, r => False), (a => 47, b => 79, p => False, o => False, r => False), (a => 111, b => 143, p => False, o => False, r => False), (a => 175, b => 207, p => False, o => False, r => False), (a => 63, b => 95, p => False, o => False, r => False), (a => 127, b => 159, p => False, o => False, r => False), (a => 191, b => 223, p => False, o => False, r => False), (a => 264, b => 272, p => False, o => False, r => False), (a => 280, b => 288, p => False, o => False, r => False), (a => 296, b => 304, p => False, o => False, r => False), (a => 312, b => 320, p => False, o => False, r => False), (a => 328, b => 336, p => False, o => False, r => False), (a => 268, b => 276, p => False, o => False, r => False), (a => 284, b => 292, p => False, o => False, r => False), (a => 300, b => 308, p => False, o => False, r => False), (a => 316, b => 324, p => False, o => False, r => False), (a => 332, b => 340, p => False, o => False, r => False), (a => 266, b => 274, p => False, o => False, r => False), (a => 282, b => 290, p => False, o => False, r => False), (a => 298, b => 306, p => False, o => False, r => False), (a => 314, b => 322, p => False, o => False, r => False), (a => 330, b => 338, p => False, o => False, r => False), (a => 270, b => 278, p => False, o => False, r => False), (a => 286, b => 294, p => False, o => False, r => False), (a => 302, b => 310, p => False, o => False, r => False), (a => 318, b => 326, p => False, o => False, r => False), (a => 334, b => 342, p => False, o => False, r => False), (a => 265, b => 273, p => False, o => False, r => False), (a => 281, b => 289, p => False, o => False, r => False), (a => 297, b => 305, p => False, o => False, r => False), (a => 313, b => 321, p => False, o => False, r => False), (a => 329, b => 337, p => False, o => False, r => False), (a => 269, b => 277, p => False, o => False, r => False), (a => 285, b => 293, p => False, o => False, r => False), (a => 301, b => 309, p => False, o => False, r => False), (a => 317, b => 325, p => False, o => False, r => False), (a => 333, b => 341, p => False, o => False, r => False), (a => 267, b => 275, p => False, o => False, r => False), (a => 283, b => 291, p => False, o => False, r => False), (a => 299, b => 307, p => False, o => False, r => False), (a => 315, b => 323, p => False, o => False, r => False), (a => 331, b => 339, p => False, o => False, r => False), (a => 271, b => 279, p => False, o => False, r => False), (a => 287, b => 295, p => False, o => False, r => False), (a => 303, b => 311, p => False, o => False, r => False), (a => 319, b => 327, p => False, o => False, r => False), (a => 335, b => 343, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 8, b => 263, p => True, o => False, r => False), (a => 9, b => 262, p => True, o => False, r => False), (a => 10, b => 261, p => True, o => False, r => False), (a => 11, b => 260, p => True, o => False, r => False), (a => 12, b => 259, p => True, o => False, r => False), (a => 13, b => 258, p => True, o => False, r => False), (a => 14, b => 257, p => True, o => False, r => False), (a => 15, b => 256, p => True, o => False, r => False), (a => 16, b => 255, p => True, o => False, r => False), (a => 17, b => 254, p => True, o => False, r => False), (a => 18, b => 253, p => True, o => False, r => False), (a => 19, b => 252, p => True, o => False, r => False), (a => 20, b => 251, p => True, o => False, r => False), (a => 21, b => 250, p => True, o => False, r => False), (a => 22, b => 249, p => True, o => False, r => False), (a => 23, b => 248, p => True, o => False, r => False), (a => 24, b => 247, p => True, o => False, r => False), (a => 25, b => 246, p => True, o => False, r => False), (a => 26, b => 245, p => True, o => False, r => False), (a => 27, b => 244, p => True, o => False, r => False), (a => 28, b => 243, p => True, o => False, r => False), (a => 29, b => 242, p => True, o => False, r => False), (a => 30, b => 241, p => True, o => False, r => False), (a => 31, b => 240, p => True, o => False, r => False), (a => 224, b => 239, p => True, o => False, r => False), (a => 225, b => 238, p => True, o => False, r => False), (a => 226, b => 237, p => True, o => False, r => False), (a => 227, b => 236, p => True, o => False, r => False), (a => 228, b => 235, p => True, o => False, r => False), (a => 229, b => 234, p => True, o => False, r => False), (a => 230, b => 233, p => True, o => False, r => False), (a => 231, b => 232, p => True, o => False, r => False)),
					((a => 16, b => 32, p => False, o => False, r => False), (a => 48, b => 64, p => False, o => False, r => False), (a => 80, b => 96, p => False, o => False, r => False), (a => 112, b => 128, p => False, o => False, r => False), (a => 144, b => 160, p => False, o => False, r => False), (a => 176, b => 192, p => False, o => False, r => False), (a => 208, b => 224, p => False, o => False, r => False), (a => 24, b => 40, p => False, o => False, r => False), (a => 56, b => 72, p => False, o => False, r => False), (a => 88, b => 104, p => False, o => False, r => False), (a => 120, b => 136, p => False, o => False, r => False), (a => 152, b => 168, p => False, o => False, r => False), (a => 184, b => 200, p => False, o => False, r => False), (a => 216, b => 232, p => False, o => False, r => False), (a => 20, b => 36, p => False, o => False, r => False), (a => 52, b => 68, p => False, o => False, r => False), (a => 84, b => 100, p => False, o => False, r => False), (a => 116, b => 132, p => False, o => False, r => False), (a => 148, b => 164, p => False, o => False, r => False), (a => 180, b => 196, p => False, o => False, r => False), (a => 212, b => 228, p => False, o => False, r => False), (a => 28, b => 44, p => False, o => False, r => False), (a => 60, b => 76, p => False, o => False, r => False), (a => 92, b => 108, p => False, o => False, r => False), (a => 124, b => 140, p => False, o => False, r => False), (a => 156, b => 172, p => False, o => False, r => False), (a => 188, b => 204, p => False, o => False, r => False), (a => 220, b => 236, p => False, o => False, r => False), (a => 18, b => 34, p => False, o => False, r => False), (a => 50, b => 66, p => False, o => False, r => False), (a => 82, b => 98, p => False, o => False, r => False), (a => 114, b => 130, p => False, o => False, r => False), (a => 146, b => 162, p => False, o => False, r => False), (a => 178, b => 194, p => False, o => False, r => False), (a => 210, b => 226, p => False, o => False, r => False), (a => 26, b => 42, p => False, o => False, r => False), (a => 58, b => 74, p => False, o => False, r => False), (a => 90, b => 106, p => False, o => False, r => False), (a => 122, b => 138, p => False, o => False, r => False), (a => 154, b => 170, p => False, o => False, r => False), (a => 186, b => 202, p => False, o => False, r => False), (a => 218, b => 234, p => False, o => False, r => False), (a => 22, b => 38, p => False, o => False, r => False), (a => 54, b => 70, p => False, o => False, r => False), (a => 86, b => 102, p => False, o => False, r => False), (a => 118, b => 134, p => False, o => False, r => False), (a => 150, b => 166, p => False, o => False, r => False), (a => 182, b => 198, p => False, o => False, r => False), (a => 214, b => 230, p => False, o => False, r => False), (a => 30, b => 46, p => False, o => False, r => False), (a => 62, b => 78, p => False, o => False, r => False), (a => 94, b => 110, p => False, o => False, r => False), (a => 126, b => 142, p => False, o => False, r => False), (a => 158, b => 174, p => False, o => False, r => False), (a => 190, b => 206, p => False, o => False, r => False), (a => 222, b => 238, p => False, o => False, r => False), (a => 17, b => 33, p => False, o => False, r => False), (a => 49, b => 65, p => False, o => False, r => False), (a => 81, b => 97, p => False, o => False, r => False), (a => 113, b => 129, p => False, o => False, r => False), (a => 145, b => 161, p => False, o => False, r => False), (a => 177, b => 193, p => False, o => False, r => False), (a => 209, b => 225, p => False, o => False, r => False), (a => 25, b => 41, p => False, o => False, r => False), (a => 57, b => 73, p => False, o => False, r => False), (a => 89, b => 105, p => False, o => False, r => False), (a => 121, b => 137, p => False, o => False, r => False), (a => 153, b => 169, p => False, o => False, r => False), (a => 185, b => 201, p => False, o => False, r => False), (a => 217, b => 233, p => False, o => False, r => False), (a => 21, b => 37, p => False, o => False, r => False), (a => 53, b => 69, p => False, o => False, r => False), (a => 85, b => 101, p => False, o => False, r => False), (a => 117, b => 133, p => False, o => False, r => False), (a => 149, b => 165, p => False, o => False, r => False), (a => 181, b => 197, p => False, o => False, r => False), (a => 213, b => 229, p => False, o => False, r => False), (a => 29, b => 45, p => False, o => False, r => False), (a => 61, b => 77, p => False, o => False, r => False), (a => 93, b => 109, p => False, o => False, r => False), (a => 125, b => 141, p => False, o => False, r => False), (a => 157, b => 173, p => False, o => False, r => False), (a => 189, b => 205, p => False, o => False, r => False), (a => 221, b => 237, p => False, o => False, r => False), (a => 19, b => 35, p => False, o => False, r => False), (a => 51, b => 67, p => False, o => False, r => False), (a => 83, b => 99, p => False, o => False, r => False), (a => 115, b => 131, p => False, o => False, r => False), (a => 147, b => 163, p => False, o => False, r => False), (a => 179, b => 195, p => False, o => False, r => False), (a => 211, b => 227, p => False, o => False, r => False), (a => 27, b => 43, p => False, o => False, r => False), (a => 59, b => 75, p => False, o => False, r => False), (a => 91, b => 107, p => False, o => False, r => False), (a => 123, b => 139, p => False, o => False, r => False), (a => 155, b => 171, p => False, o => False, r => False), (a => 187, b => 203, p => False, o => False, r => False), (a => 219, b => 235, p => False, o => False, r => False), (a => 23, b => 39, p => False, o => False, r => False), (a => 55, b => 71, p => False, o => False, r => False), (a => 87, b => 103, p => False, o => False, r => False), (a => 119, b => 135, p => False, o => False, r => False), (a => 151, b => 167, p => False, o => False, r => False), (a => 183, b => 199, p => False, o => False, r => False), (a => 215, b => 231, p => False, o => False, r => False), (a => 31, b => 47, p => False, o => False, r => False), (a => 63, b => 79, p => False, o => False, r => False), (a => 95, b => 111, p => False, o => False, r => False), (a => 127, b => 143, p => False, o => False, r => False), (a => 159, b => 175, p => False, o => False, r => False), (a => 191, b => 207, p => False, o => False, r => False), (a => 223, b => 239, p => False, o => False, r => False), (a => 260, b => 264, p => False, o => False, r => False), (a => 268, b => 272, p => False, o => False, r => False), (a => 276, b => 280, p => False, o => False, r => False), (a => 284, b => 288, p => False, o => False, r => False), (a => 292, b => 296, p => False, o => False, r => False), (a => 300, b => 304, p => False, o => False, r => False), (a => 308, b => 312, p => False, o => False, r => False), (a => 316, b => 320, p => False, o => False, r => False), (a => 324, b => 328, p => False, o => False, r => False), (a => 332, b => 336, p => False, o => False, r => False), (a => 340, b => 344, p => False, o => False, r => False), (a => 262, b => 266, p => False, o => False, r => False), (a => 270, b => 274, p => False, o => False, r => False), (a => 278, b => 282, p => False, o => False, r => False), (a => 286, b => 290, p => False, o => False, r => False), (a => 294, b => 298, p => False, o => False, r => False), (a => 302, b => 306, p => False, o => False, r => False), (a => 310, b => 314, p => False, o => False, r => False), (a => 318, b => 322, p => False, o => False, r => False), (a => 326, b => 330, p => False, o => False, r => False), (a => 334, b => 338, p => False, o => False, r => False), (a => 342, b => 346, p => False, o => False, r => False), (a => 261, b => 265, p => False, o => False, r => False), (a => 269, b => 273, p => False, o => False, r => False), (a => 277, b => 281, p => False, o => False, r => False), (a => 285, b => 289, p => False, o => False, r => False), (a => 293, b => 297, p => False, o => False, r => False), (a => 301, b => 305, p => False, o => False, r => False), (a => 309, b => 313, p => False, o => False, r => False), (a => 317, b => 321, p => False, o => False, r => False), (a => 325, b => 329, p => False, o => False, r => False), (a => 333, b => 337, p => False, o => False, r => False), (a => 341, b => 345, p => False, o => False, r => False), (a => 263, b => 267, p => False, o => False, r => False), (a => 271, b => 275, p => False, o => False, r => False), (a => 279, b => 283, p => False, o => False, r => False), (a => 287, b => 291, p => False, o => False, r => False), (a => 295, b => 299, p => False, o => False, r => False), (a => 303, b => 307, p => False, o => False, r => False), (a => 311, b => 315, p => False, o => False, r => False), (a => 319, b => 323, p => False, o => False, r => False), (a => 327, b => 331, p => False, o => False, r => False), (a => 335, b => 339, p => False, o => False, r => False), (a => 343, b => 347, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 259, p => True, o => False, r => False), (a => 5, b => 258, p => True, o => False, r => False), (a => 6, b => 257, p => True, o => False, r => False), (a => 7, b => 256, p => True, o => False, r => False), (a => 8, b => 255, p => True, o => False, r => False), (a => 9, b => 254, p => True, o => False, r => False), (a => 10, b => 253, p => True, o => False, r => False), (a => 11, b => 252, p => True, o => False, r => False), (a => 12, b => 251, p => True, o => False, r => False), (a => 13, b => 250, p => True, o => False, r => False), (a => 14, b => 249, p => True, o => False, r => False), (a => 15, b => 248, p => True, o => False, r => False), (a => 240, b => 247, p => True, o => False, r => False), (a => 241, b => 246, p => True, o => False, r => False), (a => 242, b => 245, p => True, o => False, r => False), (a => 243, b => 244, p => True, o => False, r => False)),
					((a => 8, b => 16, p => False, o => False, r => False), (a => 24, b => 32, p => False, o => False, r => False), (a => 40, b => 48, p => False, o => False, r => False), (a => 56, b => 64, p => False, o => False, r => False), (a => 72, b => 80, p => False, o => False, r => False), (a => 88, b => 96, p => False, o => False, r => False), (a => 104, b => 112, p => False, o => False, r => False), (a => 120, b => 128, p => False, o => False, r => False), (a => 136, b => 144, p => False, o => False, r => False), (a => 152, b => 160, p => False, o => False, r => False), (a => 168, b => 176, p => False, o => False, r => False), (a => 184, b => 192, p => False, o => False, r => False), (a => 200, b => 208, p => False, o => False, r => False), (a => 216, b => 224, p => False, o => False, r => False), (a => 232, b => 240, p => False, o => False, r => False), (a => 12, b => 20, p => False, o => False, r => False), (a => 28, b => 36, p => False, o => False, r => False), (a => 44, b => 52, p => False, o => False, r => False), (a => 60, b => 68, p => False, o => False, r => False), (a => 76, b => 84, p => False, o => False, r => False), (a => 92, b => 100, p => False, o => False, r => False), (a => 108, b => 116, p => False, o => False, r => False), (a => 124, b => 132, p => False, o => False, r => False), (a => 140, b => 148, p => False, o => False, r => False), (a => 156, b => 164, p => False, o => False, r => False), (a => 172, b => 180, p => False, o => False, r => False), (a => 188, b => 196, p => False, o => False, r => False), (a => 204, b => 212, p => False, o => False, r => False), (a => 220, b => 228, p => False, o => False, r => False), (a => 236, b => 244, p => False, o => False, r => False), (a => 10, b => 18, p => False, o => False, r => False), (a => 26, b => 34, p => False, o => False, r => False), (a => 42, b => 50, p => False, o => False, r => False), (a => 58, b => 66, p => False, o => False, r => False), (a => 74, b => 82, p => False, o => False, r => False), (a => 90, b => 98, p => False, o => False, r => False), (a => 106, b => 114, p => False, o => False, r => False), (a => 122, b => 130, p => False, o => False, r => False), (a => 138, b => 146, p => False, o => False, r => False), (a => 154, b => 162, p => False, o => False, r => False), (a => 170, b => 178, p => False, o => False, r => False), (a => 186, b => 194, p => False, o => False, r => False), (a => 202, b => 210, p => False, o => False, r => False), (a => 218, b => 226, p => False, o => False, r => False), (a => 234, b => 242, p => False, o => False, r => False), (a => 14, b => 22, p => False, o => False, r => False), (a => 30, b => 38, p => False, o => False, r => False), (a => 46, b => 54, p => False, o => False, r => False), (a => 62, b => 70, p => False, o => False, r => False), (a => 78, b => 86, p => False, o => False, r => False), (a => 94, b => 102, p => False, o => False, r => False), (a => 110, b => 118, p => False, o => False, r => False), (a => 126, b => 134, p => False, o => False, r => False), (a => 142, b => 150, p => False, o => False, r => False), (a => 158, b => 166, p => False, o => False, r => False), (a => 174, b => 182, p => False, o => False, r => False), (a => 190, b => 198, p => False, o => False, r => False), (a => 206, b => 214, p => False, o => False, r => False), (a => 222, b => 230, p => False, o => False, r => False), (a => 238, b => 246, p => False, o => False, r => False), (a => 9, b => 17, p => False, o => False, r => False), (a => 25, b => 33, p => False, o => False, r => False), (a => 41, b => 49, p => False, o => False, r => False), (a => 57, b => 65, p => False, o => False, r => False), (a => 73, b => 81, p => False, o => False, r => False), (a => 89, b => 97, p => False, o => False, r => False), (a => 105, b => 113, p => False, o => False, r => False), (a => 121, b => 129, p => False, o => False, r => False), (a => 137, b => 145, p => False, o => False, r => False), (a => 153, b => 161, p => False, o => False, r => False), (a => 169, b => 177, p => False, o => False, r => False), (a => 185, b => 193, p => False, o => False, r => False), (a => 201, b => 209, p => False, o => False, r => False), (a => 217, b => 225, p => False, o => False, r => False), (a => 233, b => 241, p => False, o => False, r => False), (a => 13, b => 21, p => False, o => False, r => False), (a => 29, b => 37, p => False, o => False, r => False), (a => 45, b => 53, p => False, o => False, r => False), (a => 61, b => 69, p => False, o => False, r => False), (a => 77, b => 85, p => False, o => False, r => False), (a => 93, b => 101, p => False, o => False, r => False), (a => 109, b => 117, p => False, o => False, r => False), (a => 125, b => 133, p => False, o => False, r => False), (a => 141, b => 149, p => False, o => False, r => False), (a => 157, b => 165, p => False, o => False, r => False), (a => 173, b => 181, p => False, o => False, r => False), (a => 189, b => 197, p => False, o => False, r => False), (a => 205, b => 213, p => False, o => False, r => False), (a => 221, b => 229, p => False, o => False, r => False), (a => 237, b => 245, p => False, o => False, r => False), (a => 11, b => 19, p => False, o => False, r => False), (a => 27, b => 35, p => False, o => False, r => False), (a => 43, b => 51, p => False, o => False, r => False), (a => 59, b => 67, p => False, o => False, r => False), (a => 75, b => 83, p => False, o => False, r => False), (a => 91, b => 99, p => False, o => False, r => False), (a => 107, b => 115, p => False, o => False, r => False), (a => 123, b => 131, p => False, o => False, r => False), (a => 139, b => 147, p => False, o => False, r => False), (a => 155, b => 163, p => False, o => False, r => False), (a => 171, b => 179, p => False, o => False, r => False), (a => 187, b => 195, p => False, o => False, r => False), (a => 203, b => 211, p => False, o => False, r => False), (a => 219, b => 227, p => False, o => False, r => False), (a => 235, b => 243, p => False, o => False, r => False), (a => 15, b => 23, p => False, o => False, r => False), (a => 31, b => 39, p => False, o => False, r => False), (a => 47, b => 55, p => False, o => False, r => False), (a => 63, b => 71, p => False, o => False, r => False), (a => 79, b => 87, p => False, o => False, r => False), (a => 95, b => 103, p => False, o => False, r => False), (a => 111, b => 119, p => False, o => False, r => False), (a => 127, b => 135, p => False, o => False, r => False), (a => 143, b => 151, p => False, o => False, r => False), (a => 159, b => 167, p => False, o => False, r => False), (a => 175, b => 183, p => False, o => False, r => False), (a => 191, b => 199, p => False, o => False, r => False), (a => 207, b => 215, p => False, o => False, r => False), (a => 223, b => 231, p => False, o => False, r => False), (a => 239, b => 247, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 262, b => 264, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 270, b => 272, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 278, b => 280, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 286, b => 288, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 294, b => 296, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 302, b => 304, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 310, b => 312, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 318, b => 320, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 326, b => 328, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 334, b => 336, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 342, b => 344, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 263, b => 265, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 271, b => 273, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 279, b => 281, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 287, b => 289, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 295, b => 297, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 303, b => 305, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 311, b => 313, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 319, b => 321, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 327, b => 329, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 335, b => 337, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 343, b => 345, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 257, p => True, o => False, r => False), (a => 3, b => 256, p => True, o => False, r => False), (a => 4, b => 255, p => True, o => False, r => False), (a => 5, b => 254, p => True, o => False, r => False), (a => 6, b => 253, p => True, o => False, r => False), (a => 7, b => 252, p => True, o => False, r => False), (a => 248, b => 251, p => True, o => False, r => False), (a => 249, b => 250, p => True, o => False, r => False)),
					((a => 4, b => 8, p => False, o => False, r => False), (a => 12, b => 16, p => False, o => False, r => False), (a => 20, b => 24, p => False, o => False, r => False), (a => 28, b => 32, p => False, o => False, r => False), (a => 36, b => 40, p => False, o => False, r => False), (a => 44, b => 48, p => False, o => False, r => False), (a => 52, b => 56, p => False, o => False, r => False), (a => 60, b => 64, p => False, o => False, r => False), (a => 68, b => 72, p => False, o => False, r => False), (a => 76, b => 80, p => False, o => False, r => False), (a => 84, b => 88, p => False, o => False, r => False), (a => 92, b => 96, p => False, o => False, r => False), (a => 100, b => 104, p => False, o => False, r => False), (a => 108, b => 112, p => False, o => False, r => False), (a => 116, b => 120, p => False, o => False, r => False), (a => 124, b => 128, p => False, o => False, r => False), (a => 132, b => 136, p => False, o => False, r => False), (a => 140, b => 144, p => False, o => False, r => False), (a => 148, b => 152, p => False, o => False, r => False), (a => 156, b => 160, p => False, o => False, r => False), (a => 164, b => 168, p => False, o => False, r => False), (a => 172, b => 176, p => False, o => False, r => False), (a => 180, b => 184, p => False, o => False, r => False), (a => 188, b => 192, p => False, o => False, r => False), (a => 196, b => 200, p => False, o => False, r => False), (a => 204, b => 208, p => False, o => False, r => False), (a => 212, b => 216, p => False, o => False, r => False), (a => 220, b => 224, p => False, o => False, r => False), (a => 228, b => 232, p => False, o => False, r => False), (a => 236, b => 240, p => False, o => False, r => False), (a => 244, b => 248, p => False, o => False, r => False), (a => 6, b => 10, p => False, o => False, r => False), (a => 14, b => 18, p => False, o => False, r => False), (a => 22, b => 26, p => False, o => False, r => False), (a => 30, b => 34, p => False, o => False, r => False), (a => 38, b => 42, p => False, o => False, r => False), (a => 46, b => 50, p => False, o => False, r => False), (a => 54, b => 58, p => False, o => False, r => False), (a => 62, b => 66, p => False, o => False, r => False), (a => 70, b => 74, p => False, o => False, r => False), (a => 78, b => 82, p => False, o => False, r => False), (a => 86, b => 90, p => False, o => False, r => False), (a => 94, b => 98, p => False, o => False, r => False), (a => 102, b => 106, p => False, o => False, r => False), (a => 110, b => 114, p => False, o => False, r => False), (a => 118, b => 122, p => False, o => False, r => False), (a => 126, b => 130, p => False, o => False, r => False), (a => 134, b => 138, p => False, o => False, r => False), (a => 142, b => 146, p => False, o => False, r => False), (a => 150, b => 154, p => False, o => False, r => False), (a => 158, b => 162, p => False, o => False, r => False), (a => 166, b => 170, p => False, o => False, r => False), (a => 174, b => 178, p => False, o => False, r => False), (a => 182, b => 186, p => False, o => False, r => False), (a => 190, b => 194, p => False, o => False, r => False), (a => 198, b => 202, p => False, o => False, r => False), (a => 206, b => 210, p => False, o => False, r => False), (a => 214, b => 218, p => False, o => False, r => False), (a => 222, b => 226, p => False, o => False, r => False), (a => 230, b => 234, p => False, o => False, r => False), (a => 238, b => 242, p => False, o => False, r => False), (a => 246, b => 250, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 13, b => 17, p => False, o => False, r => False), (a => 21, b => 25, p => False, o => False, r => False), (a => 29, b => 33, p => False, o => False, r => False), (a => 37, b => 41, p => False, o => False, r => False), (a => 45, b => 49, p => False, o => False, r => False), (a => 53, b => 57, p => False, o => False, r => False), (a => 61, b => 65, p => False, o => False, r => False), (a => 69, b => 73, p => False, o => False, r => False), (a => 77, b => 81, p => False, o => False, r => False), (a => 85, b => 89, p => False, o => False, r => False), (a => 93, b => 97, p => False, o => False, r => False), (a => 101, b => 105, p => False, o => False, r => False), (a => 109, b => 113, p => False, o => False, r => False), (a => 117, b => 121, p => False, o => False, r => False), (a => 125, b => 129, p => False, o => False, r => False), (a => 133, b => 137, p => False, o => False, r => False), (a => 141, b => 145, p => False, o => False, r => False), (a => 149, b => 153, p => False, o => False, r => False), (a => 157, b => 161, p => False, o => False, r => False), (a => 165, b => 169, p => False, o => False, r => False), (a => 173, b => 177, p => False, o => False, r => False), (a => 181, b => 185, p => False, o => False, r => False), (a => 189, b => 193, p => False, o => False, r => False), (a => 197, b => 201, p => False, o => False, r => False), (a => 205, b => 209, p => False, o => False, r => False), (a => 213, b => 217, p => False, o => False, r => False), (a => 221, b => 225, p => False, o => False, r => False), (a => 229, b => 233, p => False, o => False, r => False), (a => 237, b => 241, p => False, o => False, r => False), (a => 245, b => 249, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 15, b => 19, p => False, o => False, r => False), (a => 23, b => 27, p => False, o => False, r => False), (a => 31, b => 35, p => False, o => False, r => False), (a => 39, b => 43, p => False, o => False, r => False), (a => 47, b => 51, p => False, o => False, r => False), (a => 55, b => 59, p => False, o => False, r => False), (a => 63, b => 67, p => False, o => False, r => False), (a => 71, b => 75, p => False, o => False, r => False), (a => 79, b => 83, p => False, o => False, r => False), (a => 87, b => 91, p => False, o => False, r => False), (a => 95, b => 99, p => False, o => False, r => False), (a => 103, b => 107, p => False, o => False, r => False), (a => 111, b => 115, p => False, o => False, r => False), (a => 119, b => 123, p => False, o => False, r => False), (a => 127, b => 131, p => False, o => False, r => False), (a => 135, b => 139, p => False, o => False, r => False), (a => 143, b => 147, p => False, o => False, r => False), (a => 151, b => 155, p => False, o => False, r => False), (a => 159, b => 163, p => False, o => False, r => False), (a => 167, b => 171, p => False, o => False, r => False), (a => 175, b => 179, p => False, o => False, r => False), (a => 183, b => 187, p => False, o => False, r => False), (a => 191, b => 195, p => False, o => False, r => False), (a => 199, b => 203, p => False, o => False, r => False), (a => 207, b => 211, p => False, o => False, r => False), (a => 215, b => 219, p => False, o => False, r => False), (a => 223, b => 227, p => False, o => False, r => False), (a => 231, b => 235, p => False, o => False, r => False), (a => 239, b => 243, p => False, o => False, r => False), (a => 247, b => 251, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 263, b => 264, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 271, b => 272, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 279, b => 280, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 287, b => 288, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 295, b => 296, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 303, b => 304, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 311, b => 312, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 319, b => 320, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 327, b => 328, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 335, b => 336, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 343, b => 344, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 256, p => True, o => False, r => False), (a => 2, b => 255, p => True, o => False, r => False), (a => 3, b => 254, p => True, o => False, r => False), (a => 252, b => 253, p => True, o => False, r => False)),
					((a => 2, b => 4, p => False, o => False, r => False), (a => 6, b => 8, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 22, b => 24, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 30, b => 32, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 38, b => 40, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 46, b => 48, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 54, b => 56, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 62, b => 64, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 70, b => 72, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 78, b => 80, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 86, b => 88, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 94, b => 96, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 102, b => 104, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 110, b => 112, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 118, b => 120, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 126, b => 128, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 134, b => 136, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 142, b => 144, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 150, b => 152, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 158, b => 160, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 166, b => 168, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 174, b => 176, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 182, b => 184, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 190, b => 192, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 198, b => 200, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 206, b => 208, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 214, b => 216, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 222, b => 224, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 230, b => 232, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 238, b => 240, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 246, b => 248, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 23, b => 25, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 31, b => 33, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 39, b => 41, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 47, b => 49, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 55, b => 57, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 63, b => 65, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 71, b => 73, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 79, b => 81, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 87, b => 89, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 95, b => 97, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 103, b => 105, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 111, b => 113, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 119, b => 121, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 127, b => 129, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 135, b => 137, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 143, b => 145, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 151, b => 153, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 159, b => 161, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 167, b => 169, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 175, b => 177, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 183, b => 185, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 191, b => 193, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 199, b => 201, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 207, b => 209, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 215, b => 217, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 223, b => 225, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 231, b => 233, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 239, b => 241, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 247, b => 249, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 254, b => 349, p => True, o => False, r => False), (a => 255, b => 348, p => True, o => False, r => False), (a => 256, b => 347, p => True, o => False, r => False), (a => 257, b => 346, p => True, o => False, r => False), (a => 258, b => 345, p => True, o => False, r => False), (a => 259, b => 344, p => True, o => False, r => False), (a => 260, b => 343, p => True, o => False, r => False), (a => 261, b => 342, p => True, o => False, r => False), (a => 262, b => 341, p => True, o => False, r => False), (a => 263, b => 340, p => True, o => False, r => False), (a => 264, b => 339, p => True, o => False, r => False), (a => 265, b => 338, p => True, o => False, r => False), (a => 266, b => 337, p => True, o => False, r => False), (a => 267, b => 336, p => True, o => False, r => False), (a => 268, b => 335, p => True, o => False, r => False), (a => 269, b => 334, p => True, o => False, r => False), (a => 270, b => 333, p => True, o => False, r => False), (a => 271, b => 332, p => True, o => False, r => False), (a => 272, b => 331, p => True, o => False, r => False), (a => 273, b => 330, p => True, o => False, r => False), (a => 274, b => 329, p => True, o => False, r => False), (a => 275, b => 328, p => True, o => False, r => False), (a => 276, b => 327, p => True, o => False, r => False), (a => 277, b => 326, p => True, o => False, r => False), (a => 278, b => 325, p => True, o => False, r => False), (a => 279, b => 324, p => True, o => False, r => False), (a => 280, b => 323, p => True, o => False, r => False), (a => 281, b => 322, p => True, o => False, r => False), (a => 282, b => 321, p => True, o => False, r => False), (a => 283, b => 320, p => True, o => False, r => False), (a => 284, b => 319, p => True, o => False, r => False), (a => 285, b => 318, p => True, o => False, r => False), (a => 286, b => 317, p => True, o => False, r => False), (a => 287, b => 316, p => True, o => False, r => False), (a => 288, b => 315, p => True, o => False, r => False), (a => 289, b => 314, p => True, o => False, r => False), (a => 290, b => 313, p => True, o => False, r => False), (a => 291, b => 312, p => True, o => False, r => False), (a => 292, b => 311, p => True, o => False, r => False), (a => 293, b => 310, p => True, o => False, r => False), (a => 294, b => 309, p => True, o => False, r => False), (a => 295, b => 308, p => True, o => False, r => False), (a => 296, b => 307, p => True, o => False, r => False), (a => 297, b => 306, p => True, o => False, r => False), (a => 298, b => 305, p => True, o => False, r => False), (a => 299, b => 304, p => True, o => False, r => False), (a => 300, b => 303, p => True, o => False, r => False), (a => 301, b => 302, p => True, o => False, r => False)),
					((a => 1, b => 2, p => False, o => False, r => False), (a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 15, b => 16, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 23, b => 24, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 31, b => 32, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 39, b => 40, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 47, b => 48, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 55, b => 56, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 63, b => 64, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 71, b => 72, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 79, b => 80, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 87, b => 88, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 95, b => 96, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 103, b => 104, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 111, b => 112, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 119, b => 120, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 127, b => 128, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 135, b => 136, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 143, b => 144, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 151, b => 152, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 159, b => 160, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 167, b => 168, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 175, b => 176, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 183, b => 184, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 191, b => 192, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 199, b => 200, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 207, b => 208, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 215, b => 216, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 223, b => 224, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 231, b => 232, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 239, b => 240, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 247, b => 248, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 255, b => 350, p => True, o => False, r => False), (a => 256, b => 349, p => True, o => False, r => False), (a => 257, b => 348, p => True, o => False, r => False), (a => 258, b => 347, p => True, o => False, r => False), (a => 259, b => 346, p => True, o => False, r => False), (a => 260, b => 345, p => True, o => False, r => False), (a => 261, b => 344, p => True, o => False, r => False), (a => 262, b => 343, p => True, o => False, r => False), (a => 263, b => 342, p => True, o => False, r => False), (a => 264, b => 341, p => True, o => False, r => False), (a => 265, b => 340, p => True, o => False, r => False), (a => 266, b => 339, p => True, o => False, r => False), (a => 267, b => 338, p => True, o => False, r => False), (a => 268, b => 337, p => True, o => False, r => False), (a => 269, b => 336, p => True, o => False, r => False), (a => 270, b => 335, p => True, o => False, r => False), (a => 271, b => 334, p => True, o => False, r => False), (a => 272, b => 333, p => True, o => False, r => False), (a => 273, b => 332, p => True, o => False, r => False), (a => 274, b => 331, p => True, o => False, r => False), (a => 275, b => 330, p => True, o => False, r => False), (a => 276, b => 329, p => True, o => False, r => False), (a => 277, b => 328, p => True, o => False, r => False), (a => 278, b => 327, p => True, o => False, r => False), (a => 279, b => 326, p => True, o => False, r => False), (a => 280, b => 325, p => True, o => False, r => False), (a => 281, b => 324, p => True, o => False, r => False), (a => 282, b => 323, p => True, o => False, r => False), (a => 283, b => 322, p => True, o => False, r => False), (a => 284, b => 321, p => True, o => False, r => False), (a => 285, b => 320, p => True, o => False, r => False), (a => 286, b => 319, p => True, o => False, r => False), (a => 287, b => 318, p => True, o => False, r => False), (a => 288, b => 317, p => True, o => False, r => False), (a => 289, b => 316, p => True, o => False, r => False), (a => 290, b => 315, p => True, o => False, r => False), (a => 291, b => 314, p => True, o => False, r => False), (a => 292, b => 313, p => True, o => False, r => False), (a => 293, b => 312, p => True, o => False, r => False), (a => 294, b => 311, p => True, o => False, r => False), (a => 295, b => 310, p => True, o => False, r => False), (a => 296, b => 309, p => True, o => False, r => False), (a => 297, b => 308, p => True, o => False, r => False), (a => 298, b => 307, p => True, o => False, r => False), (a => 299, b => 306, p => True, o => False, r => False), (a => 300, b => 305, p => True, o => False, r => False), (a => 301, b => 304, p => True, o => False, r => False), (a => 302, b => 303, p => True, o => False, r => False)),
					((a => 128, b => 256, p => False, o => False, r => False), (a => 64, b => 320, p => False, o => False, r => False), (a => 32, b => 288, p => False, o => False, r => False), (a => 16, b => 272, p => False, o => False, r => False), (a => 80, b => 336, p => False, o => False, r => False), (a => 48, b => 304, p => False, o => False, r => False), (a => 8, b => 264, p => False, o => False, r => False), (a => 72, b => 328, p => False, o => False, r => False), (a => 40, b => 296, p => False, o => False, r => False), (a => 24, b => 280, p => False, o => False, r => False), (a => 88, b => 344, p => False, o => False, r => False), (a => 56, b => 312, p => False, o => False, r => False), (a => 4, b => 260, p => False, o => False, r => False), (a => 68, b => 324, p => False, o => False, r => False), (a => 36, b => 292, p => False, o => False, r => False), (a => 20, b => 276, p => False, o => False, r => False), (a => 84, b => 340, p => False, o => False, r => False), (a => 52, b => 308, p => False, o => False, r => False), (a => 12, b => 268, p => False, o => False, r => False), (a => 76, b => 332, p => False, o => False, r => False), (a => 44, b => 300, p => False, o => False, r => False), (a => 28, b => 284, p => False, o => False, r => False), (a => 92, b => 348, p => False, o => False, r => False), (a => 60, b => 316, p => False, o => False, r => False), (a => 2, b => 258, p => False, o => False, r => False), (a => 66, b => 322, p => False, o => False, r => False), (a => 34, b => 290, p => False, o => False, r => False), (a => 18, b => 274, p => False, o => False, r => False), (a => 82, b => 338, p => False, o => False, r => False), (a => 50, b => 306, p => False, o => False, r => False), (a => 10, b => 266, p => False, o => False, r => False), (a => 74, b => 330, p => False, o => False, r => False), (a => 42, b => 298, p => False, o => False, r => False), (a => 26, b => 282, p => False, o => False, r => False), (a => 90, b => 346, p => False, o => False, r => False), (a => 58, b => 314, p => False, o => False, r => False), (a => 6, b => 262, p => False, o => False, r => False), (a => 70, b => 326, p => False, o => False, r => False), (a => 38, b => 294, p => False, o => False, r => False), (a => 22, b => 278, p => False, o => False, r => False), (a => 86, b => 342, p => False, o => False, r => False), (a => 54, b => 310, p => False, o => False, r => False), (a => 14, b => 270, p => False, o => False, r => False), (a => 78, b => 334, p => False, o => False, r => False), (a => 46, b => 302, p => False, o => False, r => False), (a => 30, b => 286, p => False, o => False, r => False), (a => 94, b => 350, p => False, o => False, r => False), (a => 62, b => 318, p => False, o => False, r => False), (a => 1, b => 257, p => False, o => False, r => False), (a => 65, b => 321, p => False, o => False, r => False), (a => 33, b => 289, p => False, o => False, r => False), (a => 17, b => 273, p => False, o => False, r => False), (a => 81, b => 337, p => False, o => False, r => False), (a => 49, b => 305, p => False, o => False, r => False), (a => 9, b => 265, p => False, o => False, r => False), (a => 73, b => 329, p => False, o => False, r => False), (a => 41, b => 297, p => False, o => False, r => False), (a => 25, b => 281, p => False, o => False, r => False), (a => 89, b => 345, p => False, o => False, r => False), (a => 57, b => 313, p => False, o => False, r => False), (a => 5, b => 261, p => False, o => False, r => False), (a => 69, b => 325, p => False, o => False, r => False), (a => 37, b => 293, p => False, o => False, r => False), (a => 21, b => 277, p => False, o => False, r => False), (a => 85, b => 341, p => False, o => False, r => False), (a => 53, b => 309, p => False, o => False, r => False), (a => 13, b => 269, p => False, o => False, r => False), (a => 77, b => 333, p => False, o => False, r => False), (a => 45, b => 301, p => False, o => False, r => False), (a => 29, b => 285, p => False, o => False, r => False), (a => 93, b => 349, p => False, o => False, r => False), (a => 61, b => 317, p => False, o => False, r => False), (a => 3, b => 259, p => False, o => False, r => False), (a => 67, b => 323, p => False, o => False, r => False), (a => 35, b => 291, p => False, o => False, r => False), (a => 19, b => 275, p => False, o => False, r => False), (a => 83, b => 339, p => False, o => False, r => False), (a => 51, b => 307, p => False, o => False, r => False), (a => 11, b => 267, p => False, o => False, r => False), (a => 75, b => 331, p => False, o => False, r => False), (a => 43, b => 299, p => False, o => False, r => False), (a => 27, b => 283, p => False, o => False, r => False), (a => 91, b => 347, p => False, o => False, r => False), (a => 59, b => 315, p => False, o => False, r => False), (a => 7, b => 263, p => False, o => False, r => False), (a => 71, b => 327, p => False, o => False, r => False), (a => 39, b => 295, p => False, o => False, r => False), (a => 23, b => 279, p => False, o => False, r => False), (a => 87, b => 343, p => False, o => False, r => False), (a => 55, b => 311, p => False, o => False, r => False), (a => 15, b => 271, p => False, o => False, r => False), (a => 79, b => 335, p => False, o => False, r => False), (a => 47, b => 303, p => False, o => False, r => False), (a => 31, b => 287, p => False, o => False, r => False), (a => 95, b => 351, p => False, o => False, r => False), (a => 63, b => 319, p => False, o => False, r => False), (a => 0, b => 255, p => True, o => False, r => False), (a => 96, b => 254, p => True, o => False, r => False), (a => 97, b => 253, p => True, o => False, r => False), (a => 98, b => 252, p => True, o => False, r => False), (a => 99, b => 251, p => True, o => False, r => False), (a => 100, b => 250, p => True, o => False, r => False), (a => 101, b => 249, p => True, o => False, r => False), (a => 102, b => 248, p => True, o => False, r => False), (a => 103, b => 247, p => True, o => False, r => False), (a => 104, b => 246, p => True, o => False, r => False), (a => 105, b => 245, p => True, o => False, r => False), (a => 106, b => 244, p => True, o => False, r => False), (a => 107, b => 243, p => True, o => False, r => False), (a => 108, b => 242, p => True, o => False, r => False), (a => 109, b => 241, p => True, o => False, r => False), (a => 110, b => 240, p => True, o => False, r => False), (a => 111, b => 239, p => True, o => False, r => False), (a => 112, b => 238, p => True, o => False, r => False), (a => 113, b => 237, p => True, o => False, r => False), (a => 114, b => 236, p => True, o => False, r => False), (a => 115, b => 235, p => True, o => False, r => False), (a => 116, b => 234, p => True, o => False, r => False), (a => 117, b => 233, p => True, o => False, r => False), (a => 118, b => 232, p => True, o => False, r => False), (a => 119, b => 231, p => True, o => False, r => False), (a => 120, b => 230, p => True, o => False, r => False), (a => 121, b => 229, p => True, o => False, r => False), (a => 122, b => 228, p => True, o => False, r => False), (a => 123, b => 227, p => True, o => False, r => False), (a => 124, b => 226, p => True, o => False, r => False), (a => 125, b => 225, p => True, o => False, r => False), (a => 126, b => 224, p => True, o => False, r => False), (a => 127, b => 223, p => True, o => False, r => False), (a => 129, b => 222, p => True, o => False, r => False), (a => 130, b => 221, p => True, o => False, r => False), (a => 131, b => 220, p => True, o => False, r => False), (a => 132, b => 219, p => True, o => False, r => False), (a => 133, b => 218, p => True, o => False, r => False), (a => 134, b => 217, p => True, o => False, r => False), (a => 135, b => 216, p => True, o => False, r => False), (a => 136, b => 215, p => True, o => False, r => False), (a => 137, b => 214, p => True, o => False, r => False), (a => 138, b => 213, p => True, o => False, r => False), (a => 139, b => 212, p => True, o => False, r => False), (a => 140, b => 211, p => True, o => False, r => False), (a => 141, b => 210, p => True, o => False, r => False), (a => 142, b => 209, p => True, o => False, r => False), (a => 143, b => 208, p => True, o => False, r => False), (a => 144, b => 207, p => True, o => False, r => False), (a => 145, b => 206, p => True, o => False, r => False), (a => 146, b => 205, p => True, o => False, r => False), (a => 147, b => 204, p => True, o => False, r => False), (a => 148, b => 203, p => True, o => False, r => False), (a => 149, b => 202, p => True, o => False, r => False), (a => 150, b => 201, p => True, o => False, r => False), (a => 151, b => 200, p => True, o => False, r => False), (a => 152, b => 199, p => True, o => False, r => False), (a => 153, b => 198, p => True, o => False, r => False), (a => 154, b => 197, p => True, o => False, r => False), (a => 155, b => 196, p => True, o => False, r => False), (a => 156, b => 195, p => True, o => False, r => False), (a => 157, b => 194, p => True, o => False, r => False), (a => 158, b => 193, p => True, o => False, r => False), (a => 159, b => 192, p => True, o => False, r => False), (a => 160, b => 191, p => True, o => False, r => False), (a => 161, b => 190, p => True, o => False, r => False), (a => 162, b => 189, p => True, o => False, r => False), (a => 163, b => 188, p => True, o => False, r => False), (a => 164, b => 187, p => True, o => False, r => False), (a => 165, b => 186, p => True, o => False, r => False), (a => 166, b => 185, p => True, o => False, r => False), (a => 167, b => 184, p => True, o => False, r => False), (a => 168, b => 183, p => True, o => False, r => False), (a => 169, b => 182, p => True, o => False, r => False), (a => 170, b => 181, p => True, o => False, r => False), (a => 171, b => 180, p => True, o => False, r => False), (a => 172, b => 179, p => True, o => False, r => False), (a => 173, b => 178, p => True, o => False, r => False), (a => 174, b => 177, p => True, o => False, r => False), (a => 175, b => 176, p => True, o => False, r => False)),
					((a => 192, b => 320, p => False, o => False, r => False), (a => 64, b => 128, p => False, o => False, r => False), (a => 160, b => 288, p => False, o => False, r => False), (a => 144, b => 272, p => False, o => False, r => False), (a => 208, b => 336, p => False, o => False, r => False), (a => 176, b => 304, p => False, o => False, r => False), (a => 136, b => 264, p => False, o => False, r => False), (a => 200, b => 328, p => False, o => False, r => False), (a => 168, b => 296, p => False, o => False, r => False), (a => 152, b => 280, p => False, o => False, r => False), (a => 216, b => 344, p => False, o => False, r => False), (a => 184, b => 312, p => False, o => False, r => False), (a => 132, b => 260, p => False, o => False, r => False), (a => 196, b => 324, p => False, o => False, r => False), (a => 164, b => 292, p => False, o => False, r => False), (a => 148, b => 276, p => False, o => False, r => False), (a => 212, b => 340, p => False, o => False, r => False), (a => 180, b => 308, p => False, o => False, r => False), (a => 140, b => 268, p => False, o => False, r => False), (a => 204, b => 332, p => False, o => False, r => False), (a => 172, b => 300, p => False, o => False, r => False), (a => 156, b => 284, p => False, o => False, r => False), (a => 220, b => 348, p => False, o => False, r => False), (a => 188, b => 316, p => False, o => False, r => False), (a => 130, b => 258, p => False, o => False, r => False), (a => 194, b => 322, p => False, o => False, r => False), (a => 162, b => 290, p => False, o => False, r => False), (a => 146, b => 274, p => False, o => False, r => False), (a => 210, b => 338, p => False, o => False, r => False), (a => 178, b => 306, p => False, o => False, r => False), (a => 138, b => 266, p => False, o => False, r => False), (a => 202, b => 330, p => False, o => False, r => False), (a => 170, b => 298, p => False, o => False, r => False), (a => 154, b => 282, p => False, o => False, r => False), (a => 218, b => 346, p => False, o => False, r => False), (a => 186, b => 314, p => False, o => False, r => False), (a => 134, b => 262, p => False, o => False, r => False), (a => 198, b => 326, p => False, o => False, r => False), (a => 166, b => 294, p => False, o => False, r => False), (a => 150, b => 278, p => False, o => False, r => False), (a => 214, b => 342, p => False, o => False, r => False), (a => 182, b => 310, p => False, o => False, r => False), (a => 142, b => 270, p => False, o => False, r => False), (a => 206, b => 334, p => False, o => False, r => False), (a => 174, b => 302, p => False, o => False, r => False), (a => 158, b => 286, p => False, o => False, r => False), (a => 222, b => 350, p => False, o => False, r => False), (a => 190, b => 318, p => False, o => False, r => False), (a => 129, b => 257, p => False, o => False, r => False), (a => 193, b => 321, p => False, o => False, r => False), (a => 161, b => 289, p => False, o => False, r => False), (a => 145, b => 273, p => False, o => False, r => False), (a => 209, b => 337, p => False, o => False, r => False), (a => 177, b => 305, p => False, o => False, r => False), (a => 137, b => 265, p => False, o => False, r => False), (a => 201, b => 329, p => False, o => False, r => False), (a => 169, b => 297, p => False, o => False, r => False), (a => 153, b => 281, p => False, o => False, r => False), (a => 217, b => 345, p => False, o => False, r => False), (a => 185, b => 313, p => False, o => False, r => False), (a => 133, b => 261, p => False, o => False, r => False), (a => 197, b => 325, p => False, o => False, r => False), (a => 165, b => 293, p => False, o => False, r => False), (a => 149, b => 277, p => False, o => False, r => False), (a => 213, b => 341, p => False, o => False, r => False), (a => 181, b => 309, p => False, o => False, r => False), (a => 141, b => 269, p => False, o => False, r => False), (a => 205, b => 333, p => False, o => False, r => False), (a => 173, b => 301, p => False, o => False, r => False), (a => 157, b => 285, p => False, o => False, r => False), (a => 221, b => 349, p => False, o => False, r => False), (a => 189, b => 317, p => False, o => False, r => False), (a => 131, b => 259, p => False, o => False, r => False), (a => 195, b => 323, p => False, o => False, r => False), (a => 163, b => 291, p => False, o => False, r => False), (a => 147, b => 275, p => False, o => False, r => False), (a => 211, b => 339, p => False, o => False, r => False), (a => 179, b => 307, p => False, o => False, r => False), (a => 139, b => 267, p => False, o => False, r => False), (a => 203, b => 331, p => False, o => False, r => False), (a => 171, b => 299, p => False, o => False, r => False), (a => 155, b => 283, p => False, o => False, r => False), (a => 219, b => 347, p => False, o => False, r => False), (a => 187, b => 315, p => False, o => False, r => False), (a => 135, b => 263, p => False, o => False, r => False), (a => 199, b => 327, p => False, o => False, r => False), (a => 167, b => 295, p => False, o => False, r => False), (a => 151, b => 279, p => False, o => False, r => False), (a => 215, b => 343, p => False, o => False, r => False), (a => 183, b => 311, p => False, o => False, r => False), (a => 143, b => 271, p => False, o => False, r => False), (a => 207, b => 335, p => False, o => False, r => False), (a => 175, b => 303, p => False, o => False, r => False), (a => 159, b => 287, p => False, o => False, r => False), (a => 223, b => 351, p => False, o => False, r => False), (a => 191, b => 319, p => False, o => False, r => False), (a => 0, b => 256, p => True, o => False, r => False), (a => 1, b => 255, p => True, o => False, r => False), (a => 2, b => 254, p => True, o => False, r => False), (a => 3, b => 253, p => True, o => False, r => False), (a => 4, b => 252, p => True, o => False, r => False), (a => 5, b => 251, p => True, o => False, r => False), (a => 6, b => 250, p => True, o => False, r => False), (a => 7, b => 249, p => True, o => False, r => False), (a => 8, b => 248, p => True, o => False, r => False), (a => 9, b => 247, p => True, o => False, r => False), (a => 10, b => 246, p => True, o => False, r => False), (a => 11, b => 245, p => True, o => False, r => False), (a => 12, b => 244, p => True, o => False, r => False), (a => 13, b => 243, p => True, o => False, r => False), (a => 14, b => 242, p => True, o => False, r => False), (a => 15, b => 241, p => True, o => False, r => False), (a => 16, b => 240, p => True, o => False, r => False), (a => 17, b => 239, p => True, o => False, r => False), (a => 18, b => 238, p => True, o => False, r => False), (a => 19, b => 237, p => True, o => False, r => False), (a => 20, b => 236, p => True, o => False, r => False), (a => 21, b => 235, p => True, o => False, r => False), (a => 22, b => 234, p => True, o => False, r => False), (a => 23, b => 233, p => True, o => False, r => False), (a => 24, b => 232, p => True, o => False, r => False), (a => 25, b => 231, p => True, o => False, r => False), (a => 26, b => 230, p => True, o => False, r => False), (a => 27, b => 229, p => True, o => False, r => False), (a => 28, b => 228, p => True, o => False, r => False), (a => 29, b => 227, p => True, o => False, r => False), (a => 30, b => 226, p => True, o => False, r => False), (a => 31, b => 225, p => True, o => False, r => False), (a => 32, b => 224, p => True, o => False, r => False), (a => 33, b => 127, p => True, o => False, r => False), (a => 34, b => 126, p => True, o => False, r => False), (a => 35, b => 125, p => True, o => False, r => False), (a => 36, b => 124, p => True, o => False, r => False), (a => 37, b => 123, p => True, o => False, r => False), (a => 38, b => 122, p => True, o => False, r => False), (a => 39, b => 121, p => True, o => False, r => False), (a => 40, b => 120, p => True, o => False, r => False), (a => 41, b => 119, p => True, o => False, r => False), (a => 42, b => 118, p => True, o => False, r => False), (a => 43, b => 117, p => True, o => False, r => False), (a => 44, b => 116, p => True, o => False, r => False), (a => 45, b => 115, p => True, o => False, r => False), (a => 46, b => 114, p => True, o => False, r => False), (a => 47, b => 113, p => True, o => False, r => False), (a => 48, b => 112, p => True, o => False, r => False), (a => 49, b => 111, p => True, o => False, r => False), (a => 50, b => 110, p => True, o => False, r => False), (a => 51, b => 109, p => True, o => False, r => False), (a => 52, b => 108, p => True, o => False, r => False), (a => 53, b => 107, p => True, o => False, r => False), (a => 54, b => 106, p => True, o => False, r => False), (a => 55, b => 105, p => True, o => False, r => False), (a => 56, b => 104, p => True, o => False, r => False), (a => 57, b => 103, p => True, o => False, r => False), (a => 58, b => 102, p => True, o => False, r => False), (a => 59, b => 101, p => True, o => False, r => False), (a => 60, b => 100, p => True, o => False, r => False), (a => 61, b => 99, p => True, o => False, r => False), (a => 62, b => 98, p => True, o => False, r => False), (a => 63, b => 97, p => True, o => False, r => False), (a => 65, b => 96, p => True, o => False, r => False), (a => 66, b => 95, p => True, o => False, r => False), (a => 67, b => 94, p => True, o => False, r => False), (a => 68, b => 93, p => True, o => False, r => False), (a => 69, b => 92, p => True, o => False, r => False), (a => 70, b => 91, p => True, o => False, r => False), (a => 71, b => 90, p => True, o => False, r => False), (a => 72, b => 89, p => True, o => False, r => False), (a => 73, b => 88, p => True, o => False, r => False), (a => 74, b => 87, p => True, o => False, r => False), (a => 75, b => 86, p => True, o => False, r => False), (a => 76, b => 85, p => True, o => False, r => False), (a => 77, b => 84, p => True, o => False, r => False), (a => 78, b => 83, p => True, o => False, r => False), (a => 79, b => 82, p => True, o => False, r => False), (a => 80, b => 81, p => True, o => False, r => False)),
					((a => 192, b => 256, p => False, o => False, r => False), (a => 96, b => 160, p => False, o => False, r => False), (a => 224, b => 288, p => False, o => False, r => False), (a => 32, b => 64, p => False, o => False, r => False), (a => 80, b => 144, p => False, o => False, r => False), (a => 208, b => 272, p => False, o => False, r => False), (a => 112, b => 176, p => False, o => False, r => False), (a => 240, b => 304, p => False, o => False, r => False), (a => 72, b => 136, p => False, o => False, r => False), (a => 200, b => 264, p => False, o => False, r => False), (a => 104, b => 168, p => False, o => False, r => False), (a => 232, b => 296, p => False, o => False, r => False), (a => 88, b => 152, p => False, o => False, r => False), (a => 216, b => 280, p => False, o => False, r => False), (a => 120, b => 184, p => False, o => False, r => False), (a => 248, b => 312, p => False, o => False, r => False), (a => 68, b => 132, p => False, o => False, r => False), (a => 196, b => 260, p => False, o => False, r => False), (a => 100, b => 164, p => False, o => False, r => False), (a => 228, b => 292, p => False, o => False, r => False), (a => 84, b => 148, p => False, o => False, r => False), (a => 212, b => 276, p => False, o => False, r => False), (a => 116, b => 180, p => False, o => False, r => False), (a => 244, b => 308, p => False, o => False, r => False), (a => 76, b => 140, p => False, o => False, r => False), (a => 204, b => 268, p => False, o => False, r => False), (a => 108, b => 172, p => False, o => False, r => False), (a => 236, b => 300, p => False, o => False, r => False), (a => 92, b => 156, p => False, o => False, r => False), (a => 220, b => 284, p => False, o => False, r => False), (a => 124, b => 188, p => False, o => False, r => False), (a => 252, b => 316, p => False, o => False, r => False), (a => 66, b => 130, p => False, o => False, r => False), (a => 194, b => 258, p => False, o => False, r => False), (a => 98, b => 162, p => False, o => False, r => False), (a => 226, b => 290, p => False, o => False, r => False), (a => 82, b => 146, p => False, o => False, r => False), (a => 210, b => 274, p => False, o => False, r => False), (a => 114, b => 178, p => False, o => False, r => False), (a => 242, b => 306, p => False, o => False, r => False), (a => 74, b => 138, p => False, o => False, r => False), (a => 202, b => 266, p => False, o => False, r => False), (a => 106, b => 170, p => False, o => False, r => False), (a => 234, b => 298, p => False, o => False, r => False), (a => 90, b => 154, p => False, o => False, r => False), (a => 218, b => 282, p => False, o => False, r => False), (a => 122, b => 186, p => False, o => False, r => False), (a => 250, b => 314, p => False, o => False, r => False), (a => 70, b => 134, p => False, o => False, r => False), (a => 198, b => 262, p => False, o => False, r => False), (a => 102, b => 166, p => False, o => False, r => False), (a => 230, b => 294, p => False, o => False, r => False), (a => 86, b => 150, p => False, o => False, r => False), (a => 214, b => 278, p => False, o => False, r => False), (a => 118, b => 182, p => False, o => False, r => False), (a => 246, b => 310, p => False, o => False, r => False), (a => 78, b => 142, p => False, o => False, r => False), (a => 206, b => 270, p => False, o => False, r => False), (a => 110, b => 174, p => False, o => False, r => False), (a => 238, b => 302, p => False, o => False, r => False), (a => 94, b => 158, p => False, o => False, r => False), (a => 222, b => 286, p => False, o => False, r => False), (a => 126, b => 190, p => False, o => False, r => False), (a => 254, b => 318, p => False, o => False, r => False), (a => 65, b => 129, p => False, o => False, r => False), (a => 193, b => 257, p => False, o => False, r => False), (a => 97, b => 161, p => False, o => False, r => False), (a => 225, b => 289, p => False, o => False, r => False), (a => 81, b => 145, p => False, o => False, r => False), (a => 209, b => 273, p => False, o => False, r => False), (a => 113, b => 177, p => False, o => False, r => False), (a => 241, b => 305, p => False, o => False, r => False), (a => 73, b => 137, p => False, o => False, r => False), (a => 201, b => 265, p => False, o => False, r => False), (a => 105, b => 169, p => False, o => False, r => False), (a => 233, b => 297, p => False, o => False, r => False), (a => 89, b => 153, p => False, o => False, r => False), (a => 217, b => 281, p => False, o => False, r => False), (a => 121, b => 185, p => False, o => False, r => False), (a => 249, b => 313, p => False, o => False, r => False), (a => 69, b => 133, p => False, o => False, r => False), (a => 197, b => 261, p => False, o => False, r => False), (a => 101, b => 165, p => False, o => False, r => False), (a => 229, b => 293, p => False, o => False, r => False), (a => 85, b => 149, p => False, o => False, r => False), (a => 213, b => 277, p => False, o => False, r => False), (a => 117, b => 181, p => False, o => False, r => False), (a => 245, b => 309, p => False, o => False, r => False), (a => 77, b => 141, p => False, o => False, r => False), (a => 205, b => 269, p => False, o => False, r => False), (a => 109, b => 173, p => False, o => False, r => False), (a => 237, b => 301, p => False, o => False, r => False), (a => 93, b => 157, p => False, o => False, r => False), (a => 221, b => 285, p => False, o => False, r => False), (a => 125, b => 189, p => False, o => False, r => False), (a => 253, b => 317, p => False, o => False, r => False), (a => 67, b => 131, p => False, o => False, r => False), (a => 195, b => 259, p => False, o => False, r => False), (a => 99, b => 163, p => False, o => False, r => False), (a => 227, b => 291, p => False, o => False, r => False), (a => 83, b => 147, p => False, o => False, r => False), (a => 211, b => 275, p => False, o => False, r => False), (a => 115, b => 179, p => False, o => False, r => False), (a => 243, b => 307, p => False, o => False, r => False), (a => 75, b => 139, p => False, o => False, r => False), (a => 203, b => 267, p => False, o => False, r => False), (a => 107, b => 171, p => False, o => False, r => False), (a => 235, b => 299, p => False, o => False, r => False), (a => 91, b => 155, p => False, o => False, r => False), (a => 219, b => 283, p => False, o => False, r => False), (a => 123, b => 187, p => False, o => False, r => False), (a => 251, b => 315, p => False, o => False, r => False), (a => 71, b => 135, p => False, o => False, r => False), (a => 199, b => 263, p => False, o => False, r => False), (a => 103, b => 167, p => False, o => False, r => False), (a => 231, b => 295, p => False, o => False, r => False), (a => 87, b => 151, p => False, o => False, r => False), (a => 215, b => 279, p => False, o => False, r => False), (a => 119, b => 183, p => False, o => False, r => False), (a => 247, b => 311, p => False, o => False, r => False), (a => 79, b => 143, p => False, o => False, r => False), (a => 207, b => 271, p => False, o => False, r => False), (a => 111, b => 175, p => False, o => False, r => False), (a => 239, b => 303, p => False, o => False, r => False), (a => 95, b => 159, p => False, o => False, r => False), (a => 223, b => 287, p => False, o => False, r => False), (a => 127, b => 191, p => False, o => False, r => False), (a => 255, b => 319, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 8, b => 343, p => True, o => False, r => False), (a => 9, b => 342, p => True, o => False, r => False), (a => 10, b => 341, p => True, o => False, r => False), (a => 11, b => 340, p => True, o => False, r => False), (a => 12, b => 339, p => True, o => False, r => False), (a => 13, b => 338, p => True, o => False, r => False), (a => 14, b => 337, p => True, o => False, r => False), (a => 15, b => 336, p => True, o => False, r => False), (a => 16, b => 335, p => True, o => False, r => False), (a => 17, b => 334, p => True, o => False, r => False), (a => 18, b => 333, p => True, o => False, r => False), (a => 19, b => 332, p => True, o => False, r => False), (a => 20, b => 331, p => True, o => False, r => False), (a => 21, b => 330, p => True, o => False, r => False), (a => 22, b => 329, p => True, o => False, r => False), (a => 23, b => 328, p => True, o => False, r => False), (a => 24, b => 327, p => True, o => False, r => False), (a => 25, b => 326, p => True, o => False, r => False), (a => 26, b => 325, p => True, o => False, r => False), (a => 27, b => 324, p => True, o => False, r => False), (a => 28, b => 323, p => True, o => False, r => False), (a => 29, b => 322, p => True, o => False, r => False), (a => 30, b => 321, p => True, o => False, r => False), (a => 31, b => 320, p => True, o => False, r => False), (a => 33, b => 128, p => True, o => False, r => False), (a => 34, b => 63, p => True, o => False, r => False), (a => 35, b => 62, p => True, o => False, r => False), (a => 36, b => 61, p => True, o => False, r => False), (a => 37, b => 60, p => True, o => False, r => False), (a => 38, b => 59, p => True, o => False, r => False), (a => 39, b => 58, p => True, o => False, r => False), (a => 40, b => 57, p => True, o => False, r => False), (a => 41, b => 56, p => True, o => False, r => False), (a => 42, b => 55, p => True, o => False, r => False), (a => 43, b => 54, p => True, o => False, r => False), (a => 44, b => 53, p => True, o => False, r => False), (a => 45, b => 52, p => True, o => False, r => False), (a => 46, b => 51, p => True, o => False, r => False), (a => 47, b => 50, p => True, o => False, r => False), (a => 48, b => 49, p => True, o => False, r => False)),
					((a => 96, b => 128, p => False, o => False, r => False), (a => 160, b => 192, p => False, o => False, r => False), (a => 224, b => 256, p => False, o => False, r => False), (a => 288, b => 320, p => False, o => False, r => False), (a => 48, b => 80, p => False, o => False, r => False), (a => 112, b => 144, p => False, o => False, r => False), (a => 176, b => 208, p => False, o => False, r => False), (a => 240, b => 272, p => False, o => False, r => False), (a => 304, b => 336, p => False, o => False, r => False), (a => 16, b => 32, p => False, o => False, r => False), (a => 40, b => 72, p => False, o => False, r => False), (a => 104, b => 136, p => False, o => False, r => False), (a => 168, b => 200, p => False, o => False, r => False), (a => 232, b => 264, p => False, o => False, r => False), (a => 296, b => 328, p => False, o => False, r => False), (a => 56, b => 88, p => False, o => False, r => False), (a => 120, b => 152, p => False, o => False, r => False), (a => 184, b => 216, p => False, o => False, r => False), (a => 248, b => 280, p => False, o => False, r => False), (a => 312, b => 344, p => False, o => False, r => False), (a => 36, b => 68, p => False, o => False, r => False), (a => 100, b => 132, p => False, o => False, r => False), (a => 164, b => 196, p => False, o => False, r => False), (a => 228, b => 260, p => False, o => False, r => False), (a => 292, b => 324, p => False, o => False, r => False), (a => 52, b => 84, p => False, o => False, r => False), (a => 116, b => 148, p => False, o => False, r => False), (a => 180, b => 212, p => False, o => False, r => False), (a => 244, b => 276, p => False, o => False, r => False), (a => 308, b => 340, p => False, o => False, r => False), (a => 44, b => 76, p => False, o => False, r => False), (a => 108, b => 140, p => False, o => False, r => False), (a => 172, b => 204, p => False, o => False, r => False), (a => 236, b => 268, p => False, o => False, r => False), (a => 300, b => 332, p => False, o => False, r => False), (a => 60, b => 92, p => False, o => False, r => False), (a => 124, b => 156, p => False, o => False, r => False), (a => 188, b => 220, p => False, o => False, r => False), (a => 252, b => 284, p => False, o => False, r => False), (a => 316, b => 348, p => False, o => False, r => False), (a => 34, b => 66, p => False, o => False, r => False), (a => 98, b => 130, p => False, o => False, r => False), (a => 162, b => 194, p => False, o => False, r => False), (a => 226, b => 258, p => False, o => False, r => False), (a => 290, b => 322, p => False, o => False, r => False), (a => 50, b => 82, p => False, o => False, r => False), (a => 114, b => 146, p => False, o => False, r => False), (a => 178, b => 210, p => False, o => False, r => False), (a => 242, b => 274, p => False, o => False, r => False), (a => 306, b => 338, p => False, o => False, r => False), (a => 42, b => 74, p => False, o => False, r => False), (a => 106, b => 138, p => False, o => False, r => False), (a => 170, b => 202, p => False, o => False, r => False), (a => 234, b => 266, p => False, o => False, r => False), (a => 298, b => 330, p => False, o => False, r => False), (a => 58, b => 90, p => False, o => False, r => False), (a => 122, b => 154, p => False, o => False, r => False), (a => 186, b => 218, p => False, o => False, r => False), (a => 250, b => 282, p => False, o => False, r => False), (a => 314, b => 346, p => False, o => False, r => False), (a => 38, b => 70, p => False, o => False, r => False), (a => 102, b => 134, p => False, o => False, r => False), (a => 166, b => 198, p => False, o => False, r => False), (a => 230, b => 262, p => False, o => False, r => False), (a => 294, b => 326, p => False, o => False, r => False), (a => 54, b => 86, p => False, o => False, r => False), (a => 118, b => 150, p => False, o => False, r => False), (a => 182, b => 214, p => False, o => False, r => False), (a => 246, b => 278, p => False, o => False, r => False), (a => 310, b => 342, p => False, o => False, r => False), (a => 46, b => 78, p => False, o => False, r => False), (a => 110, b => 142, p => False, o => False, r => False), (a => 174, b => 206, p => False, o => False, r => False), (a => 238, b => 270, p => False, o => False, r => False), (a => 302, b => 334, p => False, o => False, r => False), (a => 62, b => 94, p => False, o => False, r => False), (a => 126, b => 158, p => False, o => False, r => False), (a => 190, b => 222, p => False, o => False, r => False), (a => 254, b => 286, p => False, o => False, r => False), (a => 318, b => 350, p => False, o => False, r => False), (a => 33, b => 65, p => False, o => False, r => False), (a => 97, b => 129, p => False, o => False, r => False), (a => 161, b => 193, p => False, o => False, r => False), (a => 225, b => 257, p => False, o => False, r => False), (a => 289, b => 321, p => False, o => False, r => False), (a => 49, b => 81, p => False, o => False, r => False), (a => 113, b => 145, p => False, o => False, r => False), (a => 177, b => 209, p => False, o => False, r => False), (a => 241, b => 273, p => False, o => False, r => False), (a => 305, b => 337, p => False, o => False, r => False), (a => 41, b => 73, p => False, o => False, r => False), (a => 105, b => 137, p => False, o => False, r => False), (a => 169, b => 201, p => False, o => False, r => False), (a => 233, b => 265, p => False, o => False, r => False), (a => 297, b => 329, p => False, o => False, r => False), (a => 57, b => 89, p => False, o => False, r => False), (a => 121, b => 153, p => False, o => False, r => False), (a => 185, b => 217, p => False, o => False, r => False), (a => 249, b => 281, p => False, o => False, r => False), (a => 313, b => 345, p => False, o => False, r => False), (a => 37, b => 69, p => False, o => False, r => False), (a => 101, b => 133, p => False, o => False, r => False), (a => 165, b => 197, p => False, o => False, r => False), (a => 229, b => 261, p => False, o => False, r => False), (a => 293, b => 325, p => False, o => False, r => False), (a => 53, b => 85, p => False, o => False, r => False), (a => 117, b => 149, p => False, o => False, r => False), (a => 181, b => 213, p => False, o => False, r => False), (a => 245, b => 277, p => False, o => False, r => False), (a => 309, b => 341, p => False, o => False, r => False), (a => 45, b => 77, p => False, o => False, r => False), (a => 109, b => 141, p => False, o => False, r => False), (a => 173, b => 205, p => False, o => False, r => False), (a => 237, b => 269, p => False, o => False, r => False), (a => 301, b => 333, p => False, o => False, r => False), (a => 61, b => 93, p => False, o => False, r => False), (a => 125, b => 157, p => False, o => False, r => False), (a => 189, b => 221, p => False, o => False, r => False), (a => 253, b => 285, p => False, o => False, r => False), (a => 317, b => 349, p => False, o => False, r => False), (a => 35, b => 67, p => False, o => False, r => False), (a => 99, b => 131, p => False, o => False, r => False), (a => 163, b => 195, p => False, o => False, r => False), (a => 227, b => 259, p => False, o => False, r => False), (a => 291, b => 323, p => False, o => False, r => False), (a => 51, b => 83, p => False, o => False, r => False), (a => 115, b => 147, p => False, o => False, r => False), (a => 179, b => 211, p => False, o => False, r => False), (a => 243, b => 275, p => False, o => False, r => False), (a => 307, b => 339, p => False, o => False, r => False), (a => 43, b => 75, p => False, o => False, r => False), (a => 107, b => 139, p => False, o => False, r => False), (a => 171, b => 203, p => False, o => False, r => False), (a => 235, b => 267, p => False, o => False, r => False), (a => 299, b => 331, p => False, o => False, r => False), (a => 59, b => 91, p => False, o => False, r => False), (a => 123, b => 155, p => False, o => False, r => False), (a => 187, b => 219, p => False, o => False, r => False), (a => 251, b => 283, p => False, o => False, r => False), (a => 315, b => 347, p => False, o => False, r => False), (a => 39, b => 71, p => False, o => False, r => False), (a => 103, b => 135, p => False, o => False, r => False), (a => 167, b => 199, p => False, o => False, r => False), (a => 231, b => 263, p => False, o => False, r => False), (a => 295, b => 327, p => False, o => False, r => False), (a => 55, b => 87, p => False, o => False, r => False), (a => 119, b => 151, p => False, o => False, r => False), (a => 183, b => 215, p => False, o => False, r => False), (a => 247, b => 279, p => False, o => False, r => False), (a => 311, b => 343, p => False, o => False, r => False), (a => 47, b => 79, p => False, o => False, r => False), (a => 111, b => 143, p => False, o => False, r => False), (a => 175, b => 207, p => False, o => False, r => False), (a => 239, b => 271, p => False, o => False, r => False), (a => 303, b => 335, p => False, o => False, r => False), (a => 63, b => 95, p => False, o => False, r => False), (a => 127, b => 159, p => False, o => False, r => False), (a => 191, b => 223, p => False, o => False, r => False), (a => 255, b => 287, p => False, o => False, r => False), (a => 319, b => 351, p => False, o => False, r => False), (a => 0, b => 64, p => True, o => False, r => False), (a => 1, b => 31, p => True, o => False, r => False), (a => 2, b => 30, p => True, o => False, r => False), (a => 3, b => 29, p => True, o => False, r => False), (a => 4, b => 28, p => True, o => False, r => False), (a => 5, b => 27, p => True, o => False, r => False), (a => 6, b => 26, p => True, o => False, r => False), (a => 7, b => 25, p => True, o => False, r => False), (a => 8, b => 24, p => True, o => False, r => False), (a => 9, b => 23, p => True, o => False, r => False), (a => 10, b => 22, p => True, o => False, r => False), (a => 11, b => 21, p => True, o => False, r => False), (a => 12, b => 20, p => True, o => False, r => False), (a => 13, b => 19, p => True, o => False, r => False), (a => 14, b => 18, p => True, o => False, r => False), (a => 15, b => 17, p => True, o => False, r => False)),
					((a => 48, b => 64, p => False, o => False, r => False), (a => 80, b => 96, p => False, o => False, r => False), (a => 112, b => 128, p => False, o => False, r => False), (a => 144, b => 160, p => False, o => False, r => False), (a => 176, b => 192, p => False, o => False, r => False), (a => 208, b => 224, p => False, o => False, r => False), (a => 240, b => 256, p => False, o => False, r => False), (a => 272, b => 288, p => False, o => False, r => False), (a => 304, b => 320, p => False, o => False, r => False), (a => 24, b => 40, p => False, o => False, r => False), (a => 56, b => 72, p => False, o => False, r => False), (a => 88, b => 104, p => False, o => False, r => False), (a => 120, b => 136, p => False, o => False, r => False), (a => 152, b => 168, p => False, o => False, r => False), (a => 184, b => 200, p => False, o => False, r => False), (a => 216, b => 232, p => False, o => False, r => False), (a => 248, b => 264, p => False, o => False, r => False), (a => 280, b => 296, p => False, o => False, r => False), (a => 312, b => 328, p => False, o => False, r => False), (a => 8, b => 16, p => False, o => False, r => False), (a => 20, b => 36, p => False, o => False, r => False), (a => 52, b => 68, p => False, o => False, r => False), (a => 84, b => 100, p => False, o => False, r => False), (a => 116, b => 132, p => False, o => False, r => False), (a => 148, b => 164, p => False, o => False, r => False), (a => 180, b => 196, p => False, o => False, r => False), (a => 212, b => 228, p => False, o => False, r => False), (a => 244, b => 260, p => False, o => False, r => False), (a => 276, b => 292, p => False, o => False, r => False), (a => 308, b => 324, p => False, o => False, r => False), (a => 28, b => 44, p => False, o => False, r => False), (a => 60, b => 76, p => False, o => False, r => False), (a => 92, b => 108, p => False, o => False, r => False), (a => 124, b => 140, p => False, o => False, r => False), (a => 156, b => 172, p => False, o => False, r => False), (a => 188, b => 204, p => False, o => False, r => False), (a => 220, b => 236, p => False, o => False, r => False), (a => 252, b => 268, p => False, o => False, r => False), (a => 284, b => 300, p => False, o => False, r => False), (a => 316, b => 332, p => False, o => False, r => False), (a => 18, b => 34, p => False, o => False, r => False), (a => 50, b => 66, p => False, o => False, r => False), (a => 82, b => 98, p => False, o => False, r => False), (a => 114, b => 130, p => False, o => False, r => False), (a => 146, b => 162, p => False, o => False, r => False), (a => 178, b => 194, p => False, o => False, r => False), (a => 210, b => 226, p => False, o => False, r => False), (a => 242, b => 258, p => False, o => False, r => False), (a => 274, b => 290, p => False, o => False, r => False), (a => 306, b => 322, p => False, o => False, r => False), (a => 26, b => 42, p => False, o => False, r => False), (a => 58, b => 74, p => False, o => False, r => False), (a => 90, b => 106, p => False, o => False, r => False), (a => 122, b => 138, p => False, o => False, r => False), (a => 154, b => 170, p => False, o => False, r => False), (a => 186, b => 202, p => False, o => False, r => False), (a => 218, b => 234, p => False, o => False, r => False), (a => 250, b => 266, p => False, o => False, r => False), (a => 282, b => 298, p => False, o => False, r => False), (a => 314, b => 330, p => False, o => False, r => False), (a => 22, b => 38, p => False, o => False, r => False), (a => 54, b => 70, p => False, o => False, r => False), (a => 86, b => 102, p => False, o => False, r => False), (a => 118, b => 134, p => False, o => False, r => False), (a => 150, b => 166, p => False, o => False, r => False), (a => 182, b => 198, p => False, o => False, r => False), (a => 214, b => 230, p => False, o => False, r => False), (a => 246, b => 262, p => False, o => False, r => False), (a => 278, b => 294, p => False, o => False, r => False), (a => 310, b => 326, p => False, o => False, r => False), (a => 30, b => 46, p => False, o => False, r => False), (a => 62, b => 78, p => False, o => False, r => False), (a => 94, b => 110, p => False, o => False, r => False), (a => 126, b => 142, p => False, o => False, r => False), (a => 158, b => 174, p => False, o => False, r => False), (a => 190, b => 206, p => False, o => False, r => False), (a => 222, b => 238, p => False, o => False, r => False), (a => 254, b => 270, p => False, o => False, r => False), (a => 286, b => 302, p => False, o => False, r => False), (a => 318, b => 334, p => False, o => False, r => False), (a => 17, b => 33, p => False, o => False, r => False), (a => 49, b => 65, p => False, o => False, r => False), (a => 81, b => 97, p => False, o => False, r => False), (a => 113, b => 129, p => False, o => False, r => False), (a => 145, b => 161, p => False, o => False, r => False), (a => 177, b => 193, p => False, o => False, r => False), (a => 209, b => 225, p => False, o => False, r => False), (a => 241, b => 257, p => False, o => False, r => False), (a => 273, b => 289, p => False, o => False, r => False), (a => 305, b => 321, p => False, o => False, r => False), (a => 25, b => 41, p => False, o => False, r => False), (a => 57, b => 73, p => False, o => False, r => False), (a => 89, b => 105, p => False, o => False, r => False), (a => 121, b => 137, p => False, o => False, r => False), (a => 153, b => 169, p => False, o => False, r => False), (a => 185, b => 201, p => False, o => False, r => False), (a => 217, b => 233, p => False, o => False, r => False), (a => 249, b => 265, p => False, o => False, r => False), (a => 281, b => 297, p => False, o => False, r => False), (a => 313, b => 329, p => False, o => False, r => False), (a => 21, b => 37, p => False, o => False, r => False), (a => 53, b => 69, p => False, o => False, r => False), (a => 85, b => 101, p => False, o => False, r => False), (a => 117, b => 133, p => False, o => False, r => False), (a => 149, b => 165, p => False, o => False, r => False), (a => 181, b => 197, p => False, o => False, r => False), (a => 213, b => 229, p => False, o => False, r => False), (a => 245, b => 261, p => False, o => False, r => False), (a => 277, b => 293, p => False, o => False, r => False), (a => 309, b => 325, p => False, o => False, r => False), (a => 29, b => 45, p => False, o => False, r => False), (a => 61, b => 77, p => False, o => False, r => False), (a => 93, b => 109, p => False, o => False, r => False), (a => 125, b => 141, p => False, o => False, r => False), (a => 157, b => 173, p => False, o => False, r => False), (a => 189, b => 205, p => False, o => False, r => False), (a => 221, b => 237, p => False, o => False, r => False), (a => 253, b => 269, p => False, o => False, r => False), (a => 285, b => 301, p => False, o => False, r => False), (a => 317, b => 333, p => False, o => False, r => False), (a => 19, b => 35, p => False, o => False, r => False), (a => 51, b => 67, p => False, o => False, r => False), (a => 83, b => 99, p => False, o => False, r => False), (a => 115, b => 131, p => False, o => False, r => False), (a => 147, b => 163, p => False, o => False, r => False), (a => 179, b => 195, p => False, o => False, r => False), (a => 211, b => 227, p => False, o => False, r => False), (a => 243, b => 259, p => False, o => False, r => False), (a => 275, b => 291, p => False, o => False, r => False), (a => 307, b => 323, p => False, o => False, r => False), (a => 27, b => 43, p => False, o => False, r => False), (a => 59, b => 75, p => False, o => False, r => False), (a => 91, b => 107, p => False, o => False, r => False), (a => 123, b => 139, p => False, o => False, r => False), (a => 155, b => 171, p => False, o => False, r => False), (a => 187, b => 203, p => False, o => False, r => False), (a => 219, b => 235, p => False, o => False, r => False), (a => 251, b => 267, p => False, o => False, r => False), (a => 283, b => 299, p => False, o => False, r => False), (a => 315, b => 331, p => False, o => False, r => False), (a => 23, b => 39, p => False, o => False, r => False), (a => 55, b => 71, p => False, o => False, r => False), (a => 87, b => 103, p => False, o => False, r => False), (a => 119, b => 135, p => False, o => False, r => False), (a => 151, b => 167, p => False, o => False, r => False), (a => 183, b => 199, p => False, o => False, r => False), (a => 215, b => 231, p => False, o => False, r => False), (a => 247, b => 263, p => False, o => False, r => False), (a => 279, b => 295, p => False, o => False, r => False), (a => 311, b => 327, p => False, o => False, r => False), (a => 31, b => 47, p => False, o => False, r => False), (a => 63, b => 79, p => False, o => False, r => False), (a => 95, b => 111, p => False, o => False, r => False), (a => 127, b => 143, p => False, o => False, r => False), (a => 159, b => 175, p => False, o => False, r => False), (a => 191, b => 207, p => False, o => False, r => False), (a => 223, b => 239, p => False, o => False, r => False), (a => 255, b => 271, p => False, o => False, r => False), (a => 287, b => 303, p => False, o => False, r => False), (a => 319, b => 335, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 4, b => 347, p => True, o => False, r => False), (a => 5, b => 346, p => True, o => False, r => False), (a => 6, b => 345, p => True, o => False, r => False), (a => 7, b => 344, p => True, o => False, r => False), (a => 9, b => 343, p => True, o => False, r => False), (a => 10, b => 342, p => True, o => False, r => False), (a => 11, b => 341, p => True, o => False, r => False), (a => 12, b => 340, p => True, o => False, r => False), (a => 13, b => 339, p => True, o => False, r => False), (a => 14, b => 338, p => True, o => False, r => False), (a => 15, b => 337, p => True, o => False, r => False), (a => 32, b => 336, p => True, o => False, r => False)),
					((a => 24, b => 32, p => False, o => False, r => False), (a => 40, b => 48, p => False, o => False, r => False), (a => 56, b => 64, p => False, o => False, r => False), (a => 72, b => 80, p => False, o => False, r => False), (a => 88, b => 96, p => False, o => False, r => False), (a => 104, b => 112, p => False, o => False, r => False), (a => 120, b => 128, p => False, o => False, r => False), (a => 136, b => 144, p => False, o => False, r => False), (a => 152, b => 160, p => False, o => False, r => False), (a => 168, b => 176, p => False, o => False, r => False), (a => 184, b => 192, p => False, o => False, r => False), (a => 200, b => 208, p => False, o => False, r => False), (a => 216, b => 224, p => False, o => False, r => False), (a => 232, b => 240, p => False, o => False, r => False), (a => 248, b => 256, p => False, o => False, r => False), (a => 264, b => 272, p => False, o => False, r => False), (a => 280, b => 288, p => False, o => False, r => False), (a => 296, b => 304, p => False, o => False, r => False), (a => 312, b => 320, p => False, o => False, r => False), (a => 328, b => 336, p => False, o => False, r => False), (a => 12, b => 20, p => False, o => False, r => False), (a => 28, b => 36, p => False, o => False, r => False), (a => 44, b => 52, p => False, o => False, r => False), (a => 60, b => 68, p => False, o => False, r => False), (a => 76, b => 84, p => False, o => False, r => False), (a => 92, b => 100, p => False, o => False, r => False), (a => 108, b => 116, p => False, o => False, r => False), (a => 124, b => 132, p => False, o => False, r => False), (a => 140, b => 148, p => False, o => False, r => False), (a => 156, b => 164, p => False, o => False, r => False), (a => 172, b => 180, p => False, o => False, r => False), (a => 188, b => 196, p => False, o => False, r => False), (a => 204, b => 212, p => False, o => False, r => False), (a => 220, b => 228, p => False, o => False, r => False), (a => 236, b => 244, p => False, o => False, r => False), (a => 252, b => 260, p => False, o => False, r => False), (a => 268, b => 276, p => False, o => False, r => False), (a => 284, b => 292, p => False, o => False, r => False), (a => 300, b => 308, p => False, o => False, r => False), (a => 316, b => 324, p => False, o => False, r => False), (a => 332, b => 340, p => False, o => False, r => False), (a => 4, b => 8, p => False, o => False, r => False), (a => 10, b => 18, p => False, o => False, r => False), (a => 26, b => 34, p => False, o => False, r => False), (a => 42, b => 50, p => False, o => False, r => False), (a => 58, b => 66, p => False, o => False, r => False), (a => 74, b => 82, p => False, o => False, r => False), (a => 90, b => 98, p => False, o => False, r => False), (a => 106, b => 114, p => False, o => False, r => False), (a => 122, b => 130, p => False, o => False, r => False), (a => 138, b => 146, p => False, o => False, r => False), (a => 154, b => 162, p => False, o => False, r => False), (a => 170, b => 178, p => False, o => False, r => False), (a => 186, b => 194, p => False, o => False, r => False), (a => 202, b => 210, p => False, o => False, r => False), (a => 218, b => 226, p => False, o => False, r => False), (a => 234, b => 242, p => False, o => False, r => False), (a => 250, b => 258, p => False, o => False, r => False), (a => 266, b => 274, p => False, o => False, r => False), (a => 282, b => 290, p => False, o => False, r => False), (a => 298, b => 306, p => False, o => False, r => False), (a => 314, b => 322, p => False, o => False, r => False), (a => 330, b => 338, p => False, o => False, r => False), (a => 14, b => 22, p => False, o => False, r => False), (a => 30, b => 38, p => False, o => False, r => False), (a => 46, b => 54, p => False, o => False, r => False), (a => 62, b => 70, p => False, o => False, r => False), (a => 78, b => 86, p => False, o => False, r => False), (a => 94, b => 102, p => False, o => False, r => False), (a => 110, b => 118, p => False, o => False, r => False), (a => 126, b => 134, p => False, o => False, r => False), (a => 142, b => 150, p => False, o => False, r => False), (a => 158, b => 166, p => False, o => False, r => False), (a => 174, b => 182, p => False, o => False, r => False), (a => 190, b => 198, p => False, o => False, r => False), (a => 206, b => 214, p => False, o => False, r => False), (a => 222, b => 230, p => False, o => False, r => False), (a => 238, b => 246, p => False, o => False, r => False), (a => 254, b => 262, p => False, o => False, r => False), (a => 270, b => 278, p => False, o => False, r => False), (a => 286, b => 294, p => False, o => False, r => False), (a => 302, b => 310, p => False, o => False, r => False), (a => 318, b => 326, p => False, o => False, r => False), (a => 334, b => 342, p => False, o => False, r => False), (a => 9, b => 17, p => False, o => False, r => False), (a => 25, b => 33, p => False, o => False, r => False), (a => 41, b => 49, p => False, o => False, r => False), (a => 57, b => 65, p => False, o => False, r => False), (a => 73, b => 81, p => False, o => False, r => False), (a => 89, b => 97, p => False, o => False, r => False), (a => 105, b => 113, p => False, o => False, r => False), (a => 121, b => 129, p => False, o => False, r => False), (a => 137, b => 145, p => False, o => False, r => False), (a => 153, b => 161, p => False, o => False, r => False), (a => 169, b => 177, p => False, o => False, r => False), (a => 185, b => 193, p => False, o => False, r => False), (a => 201, b => 209, p => False, o => False, r => False), (a => 217, b => 225, p => False, o => False, r => False), (a => 233, b => 241, p => False, o => False, r => False), (a => 249, b => 257, p => False, o => False, r => False), (a => 265, b => 273, p => False, o => False, r => False), (a => 281, b => 289, p => False, o => False, r => False), (a => 297, b => 305, p => False, o => False, r => False), (a => 313, b => 321, p => False, o => False, r => False), (a => 329, b => 337, p => False, o => False, r => False), (a => 13, b => 21, p => False, o => False, r => False), (a => 29, b => 37, p => False, o => False, r => False), (a => 45, b => 53, p => False, o => False, r => False), (a => 61, b => 69, p => False, o => False, r => False), (a => 77, b => 85, p => False, o => False, r => False), (a => 93, b => 101, p => False, o => False, r => False), (a => 109, b => 117, p => False, o => False, r => False), (a => 125, b => 133, p => False, o => False, r => False), (a => 141, b => 149, p => False, o => False, r => False), (a => 157, b => 165, p => False, o => False, r => False), (a => 173, b => 181, p => False, o => False, r => False), (a => 189, b => 197, p => False, o => False, r => False), (a => 205, b => 213, p => False, o => False, r => False), (a => 221, b => 229, p => False, o => False, r => False), (a => 237, b => 245, p => False, o => False, r => False), (a => 253, b => 261, p => False, o => False, r => False), (a => 269, b => 277, p => False, o => False, r => False), (a => 285, b => 293, p => False, o => False, r => False), (a => 301, b => 309, p => False, o => False, r => False), (a => 317, b => 325, p => False, o => False, r => False), (a => 333, b => 341, p => False, o => False, r => False), (a => 11, b => 19, p => False, o => False, r => False), (a => 27, b => 35, p => False, o => False, r => False), (a => 43, b => 51, p => False, o => False, r => False), (a => 59, b => 67, p => False, o => False, r => False), (a => 75, b => 83, p => False, o => False, r => False), (a => 91, b => 99, p => False, o => False, r => False), (a => 107, b => 115, p => False, o => False, r => False), (a => 123, b => 131, p => False, o => False, r => False), (a => 139, b => 147, p => False, o => False, r => False), (a => 155, b => 163, p => False, o => False, r => False), (a => 171, b => 179, p => False, o => False, r => False), (a => 187, b => 195, p => False, o => False, r => False), (a => 203, b => 211, p => False, o => False, r => False), (a => 219, b => 227, p => False, o => False, r => False), (a => 235, b => 243, p => False, o => False, r => False), (a => 251, b => 259, p => False, o => False, r => False), (a => 267, b => 275, p => False, o => False, r => False), (a => 283, b => 291, p => False, o => False, r => False), (a => 299, b => 307, p => False, o => False, r => False), (a => 315, b => 323, p => False, o => False, r => False), (a => 331, b => 339, p => False, o => False, r => False), (a => 15, b => 23, p => False, o => False, r => False), (a => 31, b => 39, p => False, o => False, r => False), (a => 47, b => 55, p => False, o => False, r => False), (a => 63, b => 71, p => False, o => False, r => False), (a => 79, b => 87, p => False, o => False, r => False), (a => 95, b => 103, p => False, o => False, r => False), (a => 111, b => 119, p => False, o => False, r => False), (a => 127, b => 135, p => False, o => False, r => False), (a => 143, b => 151, p => False, o => False, r => False), (a => 159, b => 167, p => False, o => False, r => False), (a => 175, b => 183, p => False, o => False, r => False), (a => 191, b => 199, p => False, o => False, r => False), (a => 207, b => 215, p => False, o => False, r => False), (a => 223, b => 231, p => False, o => False, r => False), (a => 239, b => 247, p => False, o => False, r => False), (a => 255, b => 263, p => False, o => False, r => False), (a => 271, b => 279, p => False, o => False, r => False), (a => 287, b => 295, p => False, o => False, r => False), (a => 303, b => 311, p => False, o => False, r => False), (a => 319, b => 327, p => False, o => False, r => False), (a => 335, b => 343, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 2, b => 349, p => True, o => False, r => False), (a => 3, b => 348, p => True, o => False, r => False), (a => 5, b => 347, p => True, o => False, r => False), (a => 6, b => 346, p => True, o => False, r => False), (a => 7, b => 345, p => True, o => False, r => False), (a => 16, b => 344, p => True, o => False, r => False)),
					((a => 12, b => 16, p => False, o => False, r => False), (a => 20, b => 24, p => False, o => False, r => False), (a => 28, b => 32, p => False, o => False, r => False), (a => 36, b => 40, p => False, o => False, r => False), (a => 44, b => 48, p => False, o => False, r => False), (a => 52, b => 56, p => False, o => False, r => False), (a => 60, b => 64, p => False, o => False, r => False), (a => 68, b => 72, p => False, o => False, r => False), (a => 76, b => 80, p => False, o => False, r => False), (a => 84, b => 88, p => False, o => False, r => False), (a => 92, b => 96, p => False, o => False, r => False), (a => 100, b => 104, p => False, o => False, r => False), (a => 108, b => 112, p => False, o => False, r => False), (a => 116, b => 120, p => False, o => False, r => False), (a => 124, b => 128, p => False, o => False, r => False), (a => 132, b => 136, p => False, o => False, r => False), (a => 140, b => 144, p => False, o => False, r => False), (a => 148, b => 152, p => False, o => False, r => False), (a => 156, b => 160, p => False, o => False, r => False), (a => 164, b => 168, p => False, o => False, r => False), (a => 172, b => 176, p => False, o => False, r => False), (a => 180, b => 184, p => False, o => False, r => False), (a => 188, b => 192, p => False, o => False, r => False), (a => 196, b => 200, p => False, o => False, r => False), (a => 204, b => 208, p => False, o => False, r => False), (a => 212, b => 216, p => False, o => False, r => False), (a => 220, b => 224, p => False, o => False, r => False), (a => 228, b => 232, p => False, o => False, r => False), (a => 236, b => 240, p => False, o => False, r => False), (a => 244, b => 248, p => False, o => False, r => False), (a => 252, b => 256, p => False, o => False, r => False), (a => 260, b => 264, p => False, o => False, r => False), (a => 268, b => 272, p => False, o => False, r => False), (a => 276, b => 280, p => False, o => False, r => False), (a => 284, b => 288, p => False, o => False, r => False), (a => 292, b => 296, p => False, o => False, r => False), (a => 300, b => 304, p => False, o => False, r => False), (a => 308, b => 312, p => False, o => False, r => False), (a => 316, b => 320, p => False, o => False, r => False), (a => 324, b => 328, p => False, o => False, r => False), (a => 332, b => 336, p => False, o => False, r => False), (a => 340, b => 344, p => False, o => False, r => False), (a => 6, b => 10, p => False, o => False, r => False), (a => 14, b => 18, p => False, o => False, r => False), (a => 22, b => 26, p => False, o => False, r => False), (a => 30, b => 34, p => False, o => False, r => False), (a => 38, b => 42, p => False, o => False, r => False), (a => 46, b => 50, p => False, o => False, r => False), (a => 54, b => 58, p => False, o => False, r => False), (a => 62, b => 66, p => False, o => False, r => False), (a => 70, b => 74, p => False, o => False, r => False), (a => 78, b => 82, p => False, o => False, r => False), (a => 86, b => 90, p => False, o => False, r => False), (a => 94, b => 98, p => False, o => False, r => False), (a => 102, b => 106, p => False, o => False, r => False), (a => 110, b => 114, p => False, o => False, r => False), (a => 118, b => 122, p => False, o => False, r => False), (a => 126, b => 130, p => False, o => False, r => False), (a => 134, b => 138, p => False, o => False, r => False), (a => 142, b => 146, p => False, o => False, r => False), (a => 150, b => 154, p => False, o => False, r => False), (a => 158, b => 162, p => False, o => False, r => False), (a => 166, b => 170, p => False, o => False, r => False), (a => 174, b => 178, p => False, o => False, r => False), (a => 182, b => 186, p => False, o => False, r => False), (a => 190, b => 194, p => False, o => False, r => False), (a => 198, b => 202, p => False, o => False, r => False), (a => 206, b => 210, p => False, o => False, r => False), (a => 214, b => 218, p => False, o => False, r => False), (a => 222, b => 226, p => False, o => False, r => False), (a => 230, b => 234, p => False, o => False, r => False), (a => 238, b => 242, p => False, o => False, r => False), (a => 246, b => 250, p => False, o => False, r => False), (a => 254, b => 258, p => False, o => False, r => False), (a => 262, b => 266, p => False, o => False, r => False), (a => 270, b => 274, p => False, o => False, r => False), (a => 278, b => 282, p => False, o => False, r => False), (a => 286, b => 290, p => False, o => False, r => False), (a => 294, b => 298, p => False, o => False, r => False), (a => 302, b => 306, p => False, o => False, r => False), (a => 310, b => 314, p => False, o => False, r => False), (a => 318, b => 322, p => False, o => False, r => False), (a => 326, b => 330, p => False, o => False, r => False), (a => 334, b => 338, p => False, o => False, r => False), (a => 342, b => 346, p => False, o => False, r => False), (a => 2, b => 4, p => False, o => False, r => False), (a => 5, b => 9, p => False, o => False, r => False), (a => 13, b => 17, p => False, o => False, r => False), (a => 21, b => 25, p => False, o => False, r => False), (a => 29, b => 33, p => False, o => False, r => False), (a => 37, b => 41, p => False, o => False, r => False), (a => 45, b => 49, p => False, o => False, r => False), (a => 53, b => 57, p => False, o => False, r => False), (a => 61, b => 65, p => False, o => False, r => False), (a => 69, b => 73, p => False, o => False, r => False), (a => 77, b => 81, p => False, o => False, r => False), (a => 85, b => 89, p => False, o => False, r => False), (a => 93, b => 97, p => False, o => False, r => False), (a => 101, b => 105, p => False, o => False, r => False), (a => 109, b => 113, p => False, o => False, r => False), (a => 117, b => 121, p => False, o => False, r => False), (a => 125, b => 129, p => False, o => False, r => False), (a => 133, b => 137, p => False, o => False, r => False), (a => 141, b => 145, p => False, o => False, r => False), (a => 149, b => 153, p => False, o => False, r => False), (a => 157, b => 161, p => False, o => False, r => False), (a => 165, b => 169, p => False, o => False, r => False), (a => 173, b => 177, p => False, o => False, r => False), (a => 181, b => 185, p => False, o => False, r => False), (a => 189, b => 193, p => False, o => False, r => False), (a => 197, b => 201, p => False, o => False, r => False), (a => 205, b => 209, p => False, o => False, r => False), (a => 213, b => 217, p => False, o => False, r => False), (a => 221, b => 225, p => False, o => False, r => False), (a => 229, b => 233, p => False, o => False, r => False), (a => 237, b => 241, p => False, o => False, r => False), (a => 245, b => 249, p => False, o => False, r => False), (a => 253, b => 257, p => False, o => False, r => False), (a => 261, b => 265, p => False, o => False, r => False), (a => 269, b => 273, p => False, o => False, r => False), (a => 277, b => 281, p => False, o => False, r => False), (a => 285, b => 289, p => False, o => False, r => False), (a => 293, b => 297, p => False, o => False, r => False), (a => 301, b => 305, p => False, o => False, r => False), (a => 309, b => 313, p => False, o => False, r => False), (a => 317, b => 321, p => False, o => False, r => False), (a => 325, b => 329, p => False, o => False, r => False), (a => 333, b => 337, p => False, o => False, r => False), (a => 341, b => 345, p => False, o => False, r => False), (a => 7, b => 11, p => False, o => False, r => False), (a => 15, b => 19, p => False, o => False, r => False), (a => 23, b => 27, p => False, o => False, r => False), (a => 31, b => 35, p => False, o => False, r => False), (a => 39, b => 43, p => False, o => False, r => False), (a => 47, b => 51, p => False, o => False, r => False), (a => 55, b => 59, p => False, o => False, r => False), (a => 63, b => 67, p => False, o => False, r => False), (a => 71, b => 75, p => False, o => False, r => False), (a => 79, b => 83, p => False, o => False, r => False), (a => 87, b => 91, p => False, o => False, r => False), (a => 95, b => 99, p => False, o => False, r => False), (a => 103, b => 107, p => False, o => False, r => False), (a => 111, b => 115, p => False, o => False, r => False), (a => 119, b => 123, p => False, o => False, r => False), (a => 127, b => 131, p => False, o => False, r => False), (a => 135, b => 139, p => False, o => False, r => False), (a => 143, b => 147, p => False, o => False, r => False), (a => 151, b => 155, p => False, o => False, r => False), (a => 159, b => 163, p => False, o => False, r => False), (a => 167, b => 171, p => False, o => False, r => False), (a => 175, b => 179, p => False, o => False, r => False), (a => 183, b => 187, p => False, o => False, r => False), (a => 191, b => 195, p => False, o => False, r => False), (a => 199, b => 203, p => False, o => False, r => False), (a => 207, b => 211, p => False, o => False, r => False), (a => 215, b => 219, p => False, o => False, r => False), (a => 223, b => 227, p => False, o => False, r => False), (a => 231, b => 235, p => False, o => False, r => False), (a => 239, b => 243, p => False, o => False, r => False), (a => 247, b => 251, p => False, o => False, r => False), (a => 255, b => 259, p => False, o => False, r => False), (a => 263, b => 267, p => False, o => False, r => False), (a => 271, b => 275, p => False, o => False, r => False), (a => 279, b => 283, p => False, o => False, r => False), (a => 287, b => 291, p => False, o => False, r => False), (a => 295, b => 299, p => False, o => False, r => False), (a => 303, b => 307, p => False, o => False, r => False), (a => 311, b => 315, p => False, o => False, r => False), (a => 319, b => 323, p => False, o => False, r => False), (a => 327, b => 331, p => False, o => False, r => False), (a => 335, b => 339, p => False, o => False, r => False), (a => 343, b => 347, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 350, p => True, o => False, r => False), (a => 3, b => 349, p => True, o => False, r => False), (a => 8, b => 348, p => True, o => False, r => False)),
					((a => 6, b => 8, p => False, o => False, r => False), (a => 10, b => 12, p => False, o => False, r => False), (a => 14, b => 16, p => False, o => False, r => False), (a => 18, b => 20, p => False, o => False, r => False), (a => 22, b => 24, p => False, o => False, r => False), (a => 26, b => 28, p => False, o => False, r => False), (a => 30, b => 32, p => False, o => False, r => False), (a => 34, b => 36, p => False, o => False, r => False), (a => 38, b => 40, p => False, o => False, r => False), (a => 42, b => 44, p => False, o => False, r => False), (a => 46, b => 48, p => False, o => False, r => False), (a => 50, b => 52, p => False, o => False, r => False), (a => 54, b => 56, p => False, o => False, r => False), (a => 58, b => 60, p => False, o => False, r => False), (a => 62, b => 64, p => False, o => False, r => False), (a => 66, b => 68, p => False, o => False, r => False), (a => 70, b => 72, p => False, o => False, r => False), (a => 74, b => 76, p => False, o => False, r => False), (a => 78, b => 80, p => False, o => False, r => False), (a => 82, b => 84, p => False, o => False, r => False), (a => 86, b => 88, p => False, o => False, r => False), (a => 90, b => 92, p => False, o => False, r => False), (a => 94, b => 96, p => False, o => False, r => False), (a => 98, b => 100, p => False, o => False, r => False), (a => 102, b => 104, p => False, o => False, r => False), (a => 106, b => 108, p => False, o => False, r => False), (a => 110, b => 112, p => False, o => False, r => False), (a => 114, b => 116, p => False, o => False, r => False), (a => 118, b => 120, p => False, o => False, r => False), (a => 122, b => 124, p => False, o => False, r => False), (a => 126, b => 128, p => False, o => False, r => False), (a => 130, b => 132, p => False, o => False, r => False), (a => 134, b => 136, p => False, o => False, r => False), (a => 138, b => 140, p => False, o => False, r => False), (a => 142, b => 144, p => False, o => False, r => False), (a => 146, b => 148, p => False, o => False, r => False), (a => 150, b => 152, p => False, o => False, r => False), (a => 154, b => 156, p => False, o => False, r => False), (a => 158, b => 160, p => False, o => False, r => False), (a => 162, b => 164, p => False, o => False, r => False), (a => 166, b => 168, p => False, o => False, r => False), (a => 170, b => 172, p => False, o => False, r => False), (a => 174, b => 176, p => False, o => False, r => False), (a => 178, b => 180, p => False, o => False, r => False), (a => 182, b => 184, p => False, o => False, r => False), (a => 186, b => 188, p => False, o => False, r => False), (a => 190, b => 192, p => False, o => False, r => False), (a => 194, b => 196, p => False, o => False, r => False), (a => 198, b => 200, p => False, o => False, r => False), (a => 202, b => 204, p => False, o => False, r => False), (a => 206, b => 208, p => False, o => False, r => False), (a => 210, b => 212, p => False, o => False, r => False), (a => 214, b => 216, p => False, o => False, r => False), (a => 218, b => 220, p => False, o => False, r => False), (a => 222, b => 224, p => False, o => False, r => False), (a => 226, b => 228, p => False, o => False, r => False), (a => 230, b => 232, p => False, o => False, r => False), (a => 234, b => 236, p => False, o => False, r => False), (a => 238, b => 240, p => False, o => False, r => False), (a => 242, b => 244, p => False, o => False, r => False), (a => 246, b => 248, p => False, o => False, r => False), (a => 250, b => 252, p => False, o => False, r => False), (a => 254, b => 256, p => False, o => False, r => False), (a => 258, b => 260, p => False, o => False, r => False), (a => 262, b => 264, p => False, o => False, r => False), (a => 266, b => 268, p => False, o => False, r => False), (a => 270, b => 272, p => False, o => False, r => False), (a => 274, b => 276, p => False, o => False, r => False), (a => 278, b => 280, p => False, o => False, r => False), (a => 282, b => 284, p => False, o => False, r => False), (a => 286, b => 288, p => False, o => False, r => False), (a => 290, b => 292, p => False, o => False, r => False), (a => 294, b => 296, p => False, o => False, r => False), (a => 298, b => 300, p => False, o => False, r => False), (a => 302, b => 304, p => False, o => False, r => False), (a => 306, b => 308, p => False, o => False, r => False), (a => 310, b => 312, p => False, o => False, r => False), (a => 314, b => 316, p => False, o => False, r => False), (a => 318, b => 320, p => False, o => False, r => False), (a => 322, b => 324, p => False, o => False, r => False), (a => 326, b => 328, p => False, o => False, r => False), (a => 330, b => 332, p => False, o => False, r => False), (a => 334, b => 336, p => False, o => False, r => False), (a => 338, b => 340, p => False, o => False, r => False), (a => 342, b => 344, p => False, o => False, r => False), (a => 346, b => 348, p => False, o => False, r => False), (a => 3, b => 5, p => False, o => False, r => False), (a => 7, b => 9, p => False, o => False, r => False), (a => 11, b => 13, p => False, o => False, r => False), (a => 15, b => 17, p => False, o => False, r => False), (a => 19, b => 21, p => False, o => False, r => False), (a => 23, b => 25, p => False, o => False, r => False), (a => 27, b => 29, p => False, o => False, r => False), (a => 31, b => 33, p => False, o => False, r => False), (a => 35, b => 37, p => False, o => False, r => False), (a => 39, b => 41, p => False, o => False, r => False), (a => 43, b => 45, p => False, o => False, r => False), (a => 47, b => 49, p => False, o => False, r => False), (a => 51, b => 53, p => False, o => False, r => False), (a => 55, b => 57, p => False, o => False, r => False), (a => 59, b => 61, p => False, o => False, r => False), (a => 63, b => 65, p => False, o => False, r => False), (a => 67, b => 69, p => False, o => False, r => False), (a => 71, b => 73, p => False, o => False, r => False), (a => 75, b => 77, p => False, o => False, r => False), (a => 79, b => 81, p => False, o => False, r => False), (a => 83, b => 85, p => False, o => False, r => False), (a => 87, b => 89, p => False, o => False, r => False), (a => 91, b => 93, p => False, o => False, r => False), (a => 95, b => 97, p => False, o => False, r => False), (a => 99, b => 101, p => False, o => False, r => False), (a => 103, b => 105, p => False, o => False, r => False), (a => 107, b => 109, p => False, o => False, r => False), (a => 111, b => 113, p => False, o => False, r => False), (a => 115, b => 117, p => False, o => False, r => False), (a => 119, b => 121, p => False, o => False, r => False), (a => 123, b => 125, p => False, o => False, r => False), (a => 127, b => 129, p => False, o => False, r => False), (a => 131, b => 133, p => False, o => False, r => False), (a => 135, b => 137, p => False, o => False, r => False), (a => 139, b => 141, p => False, o => False, r => False), (a => 143, b => 145, p => False, o => False, r => False), (a => 147, b => 149, p => False, o => False, r => False), (a => 151, b => 153, p => False, o => False, r => False), (a => 155, b => 157, p => False, o => False, r => False), (a => 159, b => 161, p => False, o => False, r => False), (a => 163, b => 165, p => False, o => False, r => False), (a => 167, b => 169, p => False, o => False, r => False), (a => 171, b => 173, p => False, o => False, r => False), (a => 175, b => 177, p => False, o => False, r => False), (a => 179, b => 181, p => False, o => False, r => False), (a => 183, b => 185, p => False, o => False, r => False), (a => 187, b => 189, p => False, o => False, r => False), (a => 191, b => 193, p => False, o => False, r => False), (a => 195, b => 197, p => False, o => False, r => False), (a => 199, b => 201, p => False, o => False, r => False), (a => 203, b => 205, p => False, o => False, r => False), (a => 207, b => 209, p => False, o => False, r => False), (a => 211, b => 213, p => False, o => False, r => False), (a => 215, b => 217, p => False, o => False, r => False), (a => 219, b => 221, p => False, o => False, r => False), (a => 223, b => 225, p => False, o => False, r => False), (a => 227, b => 229, p => False, o => False, r => False), (a => 231, b => 233, p => False, o => False, r => False), (a => 235, b => 237, p => False, o => False, r => False), (a => 239, b => 241, p => False, o => False, r => False), (a => 243, b => 245, p => False, o => False, r => False), (a => 247, b => 249, p => False, o => False, r => False), (a => 251, b => 253, p => False, o => False, r => False), (a => 255, b => 257, p => False, o => False, r => False), (a => 259, b => 261, p => False, o => False, r => False), (a => 263, b => 265, p => False, o => False, r => False), (a => 267, b => 269, p => False, o => False, r => False), (a => 271, b => 273, p => False, o => False, r => False), (a => 275, b => 277, p => False, o => False, r => False), (a => 279, b => 281, p => False, o => False, r => False), (a => 283, b => 285, p => False, o => False, r => False), (a => 287, b => 289, p => False, o => False, r => False), (a => 291, b => 293, p => False, o => False, r => False), (a => 295, b => 297, p => False, o => False, r => False), (a => 299, b => 301, p => False, o => False, r => False), (a => 303, b => 305, p => False, o => False, r => False), (a => 307, b => 309, p => False, o => False, r => False), (a => 311, b => 313, p => False, o => False, r => False), (a => 315, b => 317, p => False, o => False, r => False), (a => 319, b => 321, p => False, o => False, r => False), (a => 323, b => 325, p => False, o => False, r => False), (a => 327, b => 329, p => False, o => False, r => False), (a => 331, b => 333, p => False, o => False, r => False), (a => 335, b => 337, p => False, o => False, r => False), (a => 339, b => 341, p => False, o => False, r => False), (a => 343, b => 345, p => False, o => False, r => False), (a => 347, b => 349, p => False, o => False, r => False), (a => 1, b => 2, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 4, b => 350, p => True, o => False, r => False)),
					((a => 3, b => 4, p => False, o => False, r => False), (a => 5, b => 6, p => False, o => False, r => False), (a => 7, b => 8, p => False, o => False, r => False), (a => 9, b => 10, p => False, o => False, r => False), (a => 11, b => 12, p => False, o => False, r => False), (a => 13, b => 14, p => False, o => False, r => False), (a => 15, b => 16, p => False, o => False, r => False), (a => 17, b => 18, p => False, o => False, r => False), (a => 19, b => 20, p => False, o => False, r => False), (a => 21, b => 22, p => False, o => False, r => False), (a => 23, b => 24, p => False, o => False, r => False), (a => 25, b => 26, p => False, o => False, r => False), (a => 27, b => 28, p => False, o => False, r => False), (a => 29, b => 30, p => False, o => False, r => False), (a => 31, b => 32, p => False, o => False, r => False), (a => 33, b => 34, p => False, o => False, r => False), (a => 35, b => 36, p => False, o => False, r => False), (a => 37, b => 38, p => False, o => False, r => False), (a => 39, b => 40, p => False, o => False, r => False), (a => 41, b => 42, p => False, o => False, r => False), (a => 43, b => 44, p => False, o => False, r => False), (a => 45, b => 46, p => False, o => False, r => False), (a => 47, b => 48, p => False, o => False, r => False), (a => 49, b => 50, p => False, o => False, r => False), (a => 51, b => 52, p => False, o => False, r => False), (a => 53, b => 54, p => False, o => False, r => False), (a => 55, b => 56, p => False, o => False, r => False), (a => 57, b => 58, p => False, o => False, r => False), (a => 59, b => 60, p => False, o => False, r => False), (a => 61, b => 62, p => False, o => False, r => False), (a => 63, b => 64, p => False, o => False, r => False), (a => 65, b => 66, p => False, o => False, r => False), (a => 67, b => 68, p => False, o => False, r => False), (a => 69, b => 70, p => False, o => False, r => False), (a => 71, b => 72, p => False, o => False, r => False), (a => 73, b => 74, p => False, o => False, r => False), (a => 75, b => 76, p => False, o => False, r => False), (a => 77, b => 78, p => False, o => False, r => False), (a => 79, b => 80, p => False, o => False, r => False), (a => 81, b => 82, p => False, o => False, r => False), (a => 83, b => 84, p => False, o => False, r => False), (a => 85, b => 86, p => False, o => False, r => False), (a => 87, b => 88, p => False, o => False, r => False), (a => 89, b => 90, p => False, o => False, r => False), (a => 91, b => 92, p => False, o => False, r => False), (a => 93, b => 94, p => False, o => False, r => False), (a => 95, b => 96, p => False, o => False, r => False), (a => 97, b => 98, p => False, o => False, r => False), (a => 99, b => 100, p => False, o => False, r => False), (a => 101, b => 102, p => False, o => False, r => False), (a => 103, b => 104, p => False, o => False, r => False), (a => 105, b => 106, p => False, o => False, r => False), (a => 107, b => 108, p => False, o => False, r => False), (a => 109, b => 110, p => False, o => False, r => False), (a => 111, b => 112, p => False, o => False, r => False), (a => 113, b => 114, p => False, o => False, r => False), (a => 115, b => 116, p => False, o => False, r => False), (a => 117, b => 118, p => False, o => False, r => False), (a => 119, b => 120, p => False, o => False, r => False), (a => 121, b => 122, p => False, o => False, r => False), (a => 123, b => 124, p => False, o => False, r => False), (a => 125, b => 126, p => False, o => False, r => False), (a => 127, b => 128, p => False, o => False, r => False), (a => 129, b => 130, p => False, o => False, r => False), (a => 131, b => 132, p => False, o => False, r => False), (a => 133, b => 134, p => False, o => False, r => False), (a => 135, b => 136, p => False, o => False, r => False), (a => 137, b => 138, p => False, o => False, r => False), (a => 139, b => 140, p => False, o => False, r => False), (a => 141, b => 142, p => False, o => False, r => False), (a => 143, b => 144, p => False, o => False, r => False), (a => 145, b => 146, p => False, o => False, r => False), (a => 147, b => 148, p => False, o => False, r => False), (a => 149, b => 150, p => False, o => False, r => False), (a => 151, b => 152, p => False, o => False, r => False), (a => 153, b => 154, p => False, o => False, r => False), (a => 155, b => 156, p => False, o => False, r => False), (a => 157, b => 158, p => False, o => False, r => False), (a => 159, b => 160, p => False, o => False, r => False), (a => 161, b => 162, p => False, o => False, r => False), (a => 163, b => 164, p => False, o => False, r => False), (a => 165, b => 166, p => False, o => False, r => False), (a => 167, b => 168, p => False, o => False, r => False), (a => 169, b => 170, p => False, o => False, r => False), (a => 171, b => 172, p => False, o => False, r => False), (a => 173, b => 174, p => False, o => False, r => False), (a => 175, b => 176, p => False, o => False, r => False), (a => 177, b => 178, p => False, o => False, r => False), (a => 179, b => 180, p => False, o => False, r => False), (a => 181, b => 182, p => False, o => False, r => False), (a => 183, b => 184, p => False, o => False, r => False), (a => 185, b => 186, p => False, o => False, r => False), (a => 187, b => 188, p => False, o => False, r => False), (a => 189, b => 190, p => False, o => False, r => False), (a => 191, b => 192, p => False, o => False, r => False), (a => 193, b => 194, p => False, o => False, r => False), (a => 195, b => 196, p => False, o => False, r => False), (a => 197, b => 198, p => False, o => False, r => False), (a => 199, b => 200, p => False, o => False, r => False), (a => 201, b => 202, p => False, o => False, r => False), (a => 203, b => 204, p => False, o => False, r => False), (a => 205, b => 206, p => False, o => False, r => False), (a => 207, b => 208, p => False, o => False, r => False), (a => 209, b => 210, p => False, o => False, r => False), (a => 211, b => 212, p => False, o => False, r => False), (a => 213, b => 214, p => False, o => False, r => False), (a => 215, b => 216, p => False, o => False, r => False), (a => 217, b => 218, p => False, o => False, r => False), (a => 219, b => 220, p => False, o => False, r => False), (a => 221, b => 222, p => False, o => False, r => False), (a => 223, b => 224, p => False, o => False, r => False), (a => 225, b => 226, p => False, o => False, r => False), (a => 227, b => 228, p => False, o => False, r => False), (a => 229, b => 230, p => False, o => False, r => False), (a => 231, b => 232, p => False, o => False, r => False), (a => 233, b => 234, p => False, o => False, r => False), (a => 235, b => 236, p => False, o => False, r => False), (a => 237, b => 238, p => False, o => False, r => False), (a => 239, b => 240, p => False, o => False, r => False), (a => 241, b => 242, p => False, o => False, r => False), (a => 243, b => 244, p => False, o => False, r => False), (a => 245, b => 246, p => False, o => False, r => False), (a => 247, b => 248, p => False, o => False, r => False), (a => 249, b => 250, p => False, o => False, r => False), (a => 251, b => 252, p => False, o => False, r => False), (a => 253, b => 254, p => False, o => False, r => False), (a => 255, b => 256, p => False, o => False, r => False), (a => 257, b => 258, p => False, o => False, r => False), (a => 259, b => 260, p => False, o => False, r => False), (a => 261, b => 262, p => False, o => False, r => False), (a => 263, b => 264, p => False, o => False, r => False), (a => 265, b => 266, p => False, o => False, r => False), (a => 267, b => 268, p => False, o => False, r => False), (a => 269, b => 270, p => False, o => False, r => False), (a => 271, b => 272, p => False, o => False, r => False), (a => 273, b => 274, p => False, o => False, r => False), (a => 275, b => 276, p => False, o => False, r => False), (a => 277, b => 278, p => False, o => False, r => False), (a => 279, b => 280, p => False, o => False, r => False), (a => 281, b => 282, p => False, o => False, r => False), (a => 283, b => 284, p => False, o => False, r => False), (a => 285, b => 286, p => False, o => False, r => False), (a => 287, b => 288, p => False, o => False, r => False), (a => 289, b => 290, p => False, o => False, r => False), (a => 291, b => 292, p => False, o => False, r => False), (a => 293, b => 294, p => False, o => False, r => False), (a => 295, b => 296, p => False, o => False, r => False), (a => 297, b => 298, p => False, o => False, r => False), (a => 299, b => 300, p => False, o => False, r => False), (a => 301, b => 302, p => False, o => False, r => False), (a => 303, b => 304, p => False, o => False, r => False), (a => 305, b => 306, p => False, o => False, r => False), (a => 307, b => 308, p => False, o => False, r => False), (a => 309, b => 310, p => False, o => False, r => False), (a => 311, b => 312, p => False, o => False, r => False), (a => 313, b => 314, p => False, o => False, r => False), (a => 315, b => 316, p => False, o => False, r => False), (a => 317, b => 318, p => False, o => False, r => False), (a => 319, b => 320, p => False, o => False, r => False), (a => 321, b => 322, p => False, o => False, r => False), (a => 323, b => 324, p => False, o => False, r => False), (a => 325, b => 326, p => False, o => False, r => False), (a => 327, b => 328, p => False, o => False, r => False), (a => 329, b => 330, p => False, o => False, r => False), (a => 331, b => 332, p => False, o => False, r => False), (a => 333, b => 334, p => False, o => False, r => False), (a => 335, b => 336, p => False, o => False, r => False), (a => 337, b => 338, p => False, o => False, r => False), (a => 339, b => 340, p => False, o => False, r => False), (a => 341, b => 342, p => False, o => False, r => False), (a => 343, b => 344, p => False, o => False, r => False), (a => 345, b => 346, p => False, o => False, r => False), (a => 347, b => 348, p => False, o => False, r => False), (a => 349, b => 350, p => False, o => False, r => False), (a => 0, b => 351, p => True, o => False, r => False), (a => 1, b => 2, p => True, o => False, r => False))
				);

			when others => return empty_cfg;

		end case;
	end function get_cfg;

	function to_array(data : std_logic_vector; N : integer) return muon_a is
		variable muon : muon_a(0 to N - 1);
	begin
		for i in muon'range loop
			muon(i).pt  := data((i + 1) * word_w - 1 - IDX_WIDTH downto i * word_w);
			muon(i).idx := data((i + 1) * word_w - 1 downto i * word_w + PT_WIDTH);
		end loop;
		return muon;
	end to_array;

	function to_stdv(muon : muon_a; N : integer) return std_logic_vector is
		variable vector : std_logic_vector(N * word_w - 1 downto 0);
	begin
		for i in muon'range loop
			vector((i + 1) * word_w - 1 - IDX_WIDTH downto i * word_w) := muon(i).pt;
			vector((i + 1) * word_w - 1 downto i * word_w + PT_WIDTH)  := muon(i).idx;
		end loop;
		return vector;
	end to_stdv;

end package body csn_pkg;
